`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hRa0GRImT8YcQlmWFV+vMHYSsEI52cyMWmcxzY6IAm+ZyXJNrpxT0ixlgWDJ/EgFAY2YhIam/tzK
N9c4uoFk7A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZIZn6elsuGvDqXXgH+2znh/3m25gw8eMgiW6h/D2XAX8pAbVOqTpaaAu8lyhmwCNkRMAhEVzIjUT
0v67Hn2IAnoNrsGSjcYowIw8WPquzBC0O32To+o2XQDesiPm2n0EA33VJ5HOOKNC9eVIs7b90yaN
BlgWT58+XJuLuhSniV4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FC6THI0G35SGPQEJh9JkbUmH5FoUwqOxzexRACJ39PALi3OmCgBmGl9nRsKp98Zhv6S6lRJi5m+U
oa1FxJiZCC2t7O1GPEIJgmPLY/PbYoiMs0BSfwLEGso5HEaEDtKYzOxVlMeduP8O1vGu6XRvduWO
L8Xrgsu6cFKn9Oz4TvyMy8fS4BKOOMIYHk+AvE4WUr4ZPwI9g0pw0NzIkFHnh/59YB1IdRI6dcHn
A69IWI/zBtD9hvDC3buv1d7YXfZGLYXj1zcWgE5iFw3OANIJ/3wwoY/G9Spe1quwZAX7qEVOw7j4
ey/SXS49JmXfcL6TXyb4+T6zbrjGPHAyYJwRIg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PBxjocOlJwBpwIFDR28jk7BESYWFC6ML1qwzlwrw6V48UFZGXGe3d7xjmMwsRYRIUXCtO+CB6BfD
BuDWw0llGpVhWp4gxCzi77C3X4JyuWxkaoQeqSKfPnx4d2rr+v0YO5DZqNZFCjySSD3drVL1sPjC
dX5PrpB1gemAkEF9DpSK2Pz14H8OyMZ7ysIpZGPwN7b+K6v356waWSK6A9cQZgwvZbNsby1Ypgzy
bVMA1m7yCr24wfHxY1bPiGFIr8ikzSu6IrnxwSWcRhJXBjMuQvK91C7i3JwAUzBQMJlP91ApQdAF
/HktGGZXkzE1ZAFwfG7VG9gmvJko2oEyRYIZow==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
D3iiskMSAmhggSdSRKuuAs7X55v9whKqZ3poDY4/UVjilEIhk0AZPl9Go1ErgGkier6QCJvoo7uW
s1JCbXuZRPjqFovsugIQjVHP6DcT8K57QMEwdHu2ybXpP/Lmhgg13n+UeQWQzlkK0WOcvXLEOT0k
3lh6qo8OsHtm0IiN5X631AQ96O5CdVJuU4fd/S9cZjPFRhoWbvKViTdVSJOfTD+LCCaR27xZCsE7
7irfraBbSY3/g748jREDJDl8dg3s39OMQECe1Gc/eO87dmMHyOUSMREIRHgIDnFz61l1ctPIvPcr
yrarHfOF07k4wO/3Sf1Ezu43mRFkVA7+J5M8Mg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VY11L2vkFT3Fqdzmb5pPrvvcekipOFwuApdkldlZDTmW4ugweAD3PnxqNh6dGtjLHBrjVjv1Mdfy
Xikp9dY0NuHQGrriGlFvnC8Qs9saTcduZXB5+v2+NabX6MIAp8gEOmS2z2sNuX6C6HhC+X97Avvi
Sfs6Dazhq5mXriaXI4U=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
H4r0uFGQA1yIbVPIb59MnCh++12qcAESGLrt0S24zf4znjh0AzrJlyVnkhrA7mxT6iHKi0NgFFMA
W4K0W+wYysidfkmvYZenPHZSDPuHt6mv1pF4SJ645ug3mBxdGB2h4D/Zzn9aLso4TOca4QOLW32j
RLj1cXkpF8oD//8wKzMYORTjKiDttvnl5W6jOfIXPxo7VbrAOsVpsFXlFKn/G0ptiLHVEu0U/Vxl
yaKsYOQsNXSw3RiONZ+cflAm5BOea1rmTNS69lo++pjQAfkYwDXr1M1hoYjteEVfg9DaK8OSRMyE
Y4jk3H3OpztNRmMbUbGFdU9Qjtfh0bh2lamnWw==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DHMpgf3HyOeA2ZRozTpXOZcMkD7fDghjVjp9qR/joma/4HuQpBqINHeUc5wSaoK2ocniM4fX48dr
4NV8hPskDDZp7+c88GxnQmdbzfv6O6e9PbKbYpdkBkj/gzmJc2CZtdMuc9QQHdv3bWDKNuGAlQAD
LIZTzm2Exj1vAgLBf/olc7ekW0p/Vq3QdFAiR6A8fGrCrd+UEcCoydkzOmn7JSAxiYOKdjs0xJ2T
FhvbzExS3UIyghTUHVx6dXpETh26W1xRKwYTVz0GZehUrHEKrYU7WiD899nLcAgVAHXHkxjcIPkx
TEntACr92IGrhqpicKLyonsGYS3JhiXAYdTcxg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 859744)
`protect data_block
ZnTBxNa08UepqAz19wcl78ScRlPB7vYHWF47S3PukMDXIKFR4u+RV8THSuSgl/mRgphtRNH62cE2
DlANHNA2oKzzopOduzu+N9FVs1/xK1k3pzl1mwzIseKPMAyHFc6UOENcvjio3ZvBRPauP45Sd3N9
j6EZ9jXn9als3G9Ry0NnCkdbIWst/3Z0QtjGjtaPcLoQw860vFCcFxBvKMnjQVFUWY4HDv+1MeJD
oxTuGYitbKuzH6GiXRDasbTEfztQZHp0+gleYEk3+xMFYaNWZySG9s2MLCzrI3Af5YKS80zHYHmV
w4wEletjzrmRQeJ/8eicqvAvN30AxIG3qkAIGcvHRySe5Xc6DtLv0qZmo+5J0jitVtoe1i1T4F+d
IquET6BLl5hg+1tmp1/uoS3tFsOPZhsW1LFOubNoZa/epdp4PlnNR9R1R6s6Ms++K9zBtP7xOzXj
/Qe6tfasGZHBTQCX9Wh86sRaPh5IKs9fyUBx2Re6XHqxLeIk3YhUAbsGuzdOUX6E1JfAS4qzum4x
J4aYcGJkDNixNa7r9HpQf82zpU3FwzsG59q38IknFU80iDvZuBoq8VmGQRmdzXE1poK+hpq84l9B
Y97YvugnES/hli6j6fnvgrg9LWPgehT4W2GRz36EV9IQ3QTmUdcuR6PmYpeVYfVKz0tv079uW4MG
FKBZDeBgTj/EuVh8u3WMBFQ0PcMr45MuzdPpOdRnts9UmcFj6yDBNwXO0YlBrIYNK6r7mAdKUioW
svxFHnbMRElLHiRa1fV/ia/YnKk0M+uKZ3JXFQWv1OjT/pCzpvChK5fnbUglnwzL/q2D3kPAkzKL
U9UuAVH9Dmnb2CKT4KjVyA0ifDQcWM+KM/51qWvVSlkw+aKgybegS/KGK/i/yUpJHeIMGd3X5UaC
CmUgRaNYhTA/vYkds4xYlczJlsAUjtZx4WdDTvVuuxSnFuRO2YRTp4Lz5cgBU9YhM9JHLliWvdJD
sfF23SId+wBonBquWFXT+RzeCRs/lpz3qzhZeGvs5HlfDpSPYGoDup3nvKUwN3oznB3E+rtzc7RH
M8ePlw60LfkIdc0x4HaaPC6P0+JY7GjPHwtvERcbBoBa087HIsZtK+zO2onLcEpdsOTxAZXMeHOi
AWfoub5kAXA9CsqDROraBFRV7DZQQibMyE47cQrLaJ+qct/aCZRVazfoFNDXjaSZzKxxBELe8bUv
935huJ5FrplkCoNC2YBun/RpAfC1cADIWKVdfOpZWnx5a9BGLl2nOJcxCkwekuCOlpEfhNrNdKHa
xKOb9xe2PhwKvrTurD27nE7Z1guc5aMlJipv7S7FBpdWU0FND4jiLIktygZkypGaEYe73r5TnWuE
r1lhMBnl6nE8ndR9QoKXwb10Pw20JnD717CCvLvbMBaU8tjxhK5467y2nmLr2dADv1dLmDg7G3t8
tWV2DShRiF1XutDRn3kLZwqMbFroTnd1Ib6XImQnUew6WRKhiwjySJvqceNrpW63+Dt5cA4eDeF1
QBN5Or0UmT0Kfyj38tuwXgP7YbOvzLFAon1A3e9hvHdKHxcYYb/Jo2EopdzN3klWaTY1OIXgvrhO
1yMDhhBh8wLWTCRRQncb5Mkvmx11tDCwh2+L//YbhS1kE34g/9HbvB//HHQg9zBcJnW7T0rFv7L7
LdJC1YextxnDlnbMCsYzAl1DbGJzY0/qvAz9+mz210rcGEj6SP8sNblPjH99WmxUBnzwmjLh5uJg
Z2+8iklglDTHFPGkljoVmS/LgG5e+HiOJ838jJlGAX0+FHAiuTn1WvH5iTSeLHRWkRAqCzEM3tAZ
JkqI+kI2EW7U223QFF0VH/sVHXwMdb1hjZUFI7k4sVvd9CP6EQm3rTcSSLFCMRy8mMBlukvJwQTu
cSRN52t+wIWO4/YhYOhnmapZg9xW/tqsRAE3MQfEnFWs82B8lGBWW/fE+yIFs4KoMDOrlueJHtij
LdvCHh00flgl39QdXwYeYVFrs91VvhdEhScAM0Fo6RwhJ11AqveKoNEz25Bj+uIjQuqmhIawDY9T
Ha5Ax7jxnwn7nD2M0DPDFQDVLvem9rY33a1N8ivxq/i6tuo0qRzBFUD51nMZwDIW8jzNqeiff4R0
QD+bVJfaDfcZ9O3nzZ2DP4qY8WqXx0ElIvBOtzbmsUZYbEBCLYNuTHRzLNBqMnPmH4nerM8kt3IC
DO/rjmJ2w/DgbbYnI/N5iK8Lz6Lt+FZdayRxgb261ywq4JG0q1sMYZOxGtV24PfusNW6w0pgHh45
Ytrzmc02vTbi1rLa4QVbASq7KGLx9wzuh+maX9tGmyoB56SCQiSIiZqdJQ9/osQ/GckIHS1wGy14
jeRvNR2kUzffkAeLzUw3L7n9k7kg06lW44HNetRsHIEY3Q7pbfKAjHxbVyrM9MKhUQY8bsUazN8q
WRiCVFQOZjr0gsaQV4PPnz4vsroNR+8OUyi7/crCNenUNQAlcaz3+Zse+BsNK2LCxVD83sTsOlkl
i5kGtfrDjQQBXnUj03ui5x1Ft8T9XoGyCS0VbMKhq5mY/qU38tHffbyy6OHDlxuxqudOxmpYzT1/
+3GhpZgJ/rowok2Bc9vyWfGb8L+86rERrjTSjDKth1i9HJ1Vi+Fabr6UliK85zK/Lgv/UXjjeF8O
9rsBUNvii0nAOYe4h6uzJwZsJ7WY6OQLtsa/Q9HnjEi8kP3llIaDQ+m9uUZIRfw/BZImk3g8Djl0
dySEnsNqQuRtiZwsCy91HQL3lq+7BAmRxFBWCMbn8+5IjceDtbokklnE3HYEBWGuuQ1R2kDccuG/
KMUSlwpHOUfYMrdDZPJepH1hUFSKh8E4gpVVVGMWIY0KcRE6nytrZ+smJFn86c2po9vqeVNbacjp
xoPgIUoBJzWIJxAC+TD0HB0bJYhsG/Wqdr6ROc4O47sBe7AhMxUYBfARynqw9kjW1h2FII6ZgrNa
zEOjHzwx+1gt3SN0d61RMmWjFpaZoPUJExuCushhd3E3OGtC9aiSfxQwt1AOSv5aywr6nAc2lvBp
06O5JVV9w5mCyrfjKzvjBaZ4jfHZxcFnGldFSWOQElrMlFRapBnn5X/gEuKN3V3s1tKXwPQdg9mA
4zDQmpV7RfsOPwrubRDet3kh993TTpz7eFR9z0gLrCcYarXpL8e29e6IhbSMv/9dU0CVALsKdHlE
Rrc+LHYXx2F0LDL80UMS218nN/Hab9dY8SXXCCwU41Juu+fO9UwIat/u06nsWdnvAab30bwnWysL
uykVln1yLwAT/fuafvOVVS7zdH+rrO8+fGUdi48DG+AUT4NKyG7AkN1KEen2HmH8A4dEN102G8EU
9jRRoCSW6L5a/X8sFSm0XkMxSgJ1rZNKCzDYs/fr5aEvu8Qn8VNBivn5+dAJYsLkmaeGZKxBpe2G
Zm9cuDN8a6xAGa5PdNoiPOTC4ECm4XkiZUgUuakbvDn255fIn4iM+7xmpzxj5M7H8COn5xBvuaHK
1acJmWJVl9bb0VINctxuABiLVoqc42Y8gDWrM1u49lpzbB3uK2DYH+7SKrkKj0LBckIduVoiTQhs
FUq9Zo9UQ8vQWKCtpQ11Z63o3W6t5+yWM4JNPhdGVqO1Mdprjc416ajD56z+QpSdpiFo1uNN02QP
f45wWYfDjLPNL6i94+z7HfiY9v1LvkzZliwj45o9Y8Ez7PX5da5GmpgxooEk6GFVToEMlLEebGrI
NdfJ3e1MeGnwnKeSEKblnGJO/SHGULi5xWX9fi2oIzcRrF17r3SeUeEELEwe+qCsumFLXdRoPP0a
p3gGr8c93nvhnYDHKx3d1+fqwaPbgDUCFYdswF6ydguLaPbbonHlGpQhqhQUQOTVzylHj3WluDc8
7oqHo1VT+d0PpSEPzfFiOIIN3XzSObo4F7yUbgBGNJpHehlntru7BCFXBCSzWocmgS+ufqrRkN2g
QTL8dqhUw4IvqCJKbebSgWTi6j7OocWLYB6/jcT4dvNtXPqkccTNq/Jd5DHqOYdgfjaED3vSgDSN
z/FjogZTYKt+lPs4rW2XaeIbFmnEdW7CCdDNORoJdMkjGvzNj6ikyzAKMwSGVZY9h+7LXSlIX/Zm
Ei6hsLv/5pUQS0zSFgjLAD/0dJLy6OZvSys0zFcr2OqtXYFclQ4UeNjoFLm6Yn464sTstR/mBNao
fYeJsgHzL1liWBYw9MV5c959PxNHL2nHcPdiSOiw8ZyTVNrrj5HgMuGIRqIYU6r3ePYS5m1MzF3T
Kpqx29n97hJ46aOhMwHrJovMJuZSIVUu4a4m2xwx3OAfCo345ZHCOQLM21vfisIWyRzp30JOO3mM
woyqMrWEJFSgTprsJMqgkT7VUVwoaKWU8rGDiNuLUyiT6rxixE/N+YcwARp7DYbT+rte2F4M/b4W
xon6N+C5HaXF7IpsJcaBnirkTg9L5ngwkwVdpt7CKwl90D56bvKrhk0oNW+UyQfcSz8swgFOYRYE
1CpvSFXgQtHapq/raZj9kAyB0lB/BnVNoMFzMFwI5xW0hi/CZHws8Aj+uVXwYmuREKz+5sOlvqE/
TeiUDT23FnZ8CTLklzAam5KpW/AqDi7sKI18E4BF0XQ+QH89a2XrYH6S5jJFFY7BZzrCrWxW+0xI
F1LLbIw3I0Adc79NJQHcCSsWGwAVVEiHzTTsKYNgEetj97n1aUMgKdeKX/E+tYC4zGRHFkIDAhSv
K8OFn8U+lT7HDETQYpTHFKc9xHALQUiEEfIb+iAVpharkrf2v7dO4+fJOoFVT1sdQedxmpLoV2v4
wYCPizD16nPaWxeqJnyF1ORRirIdVaCt8m5Lxr/GVas5w1AtCZBAmcTCqMIOg+g86CTy9wh2iAGL
eVTfpE1ktRN8ghxVJaYFui+taD9JTaySR462s3v9UOep1uC0hFSWFk0osUBFBIY9jOXnS0C2PZyB
sQpRkkolW2qMtJGh9BkvazsVt2dgGjHdz3e4ZMYehTYatKJpE6zCJ3pj2cD/s8/lf9jsZchhzJ3B
4ncMrN0TUsBai/mTrkwkPkOS2V40FVAKta7FmdJQmQOcXMU7i1tSCrfbKWohu9Xg23YnQcrm4Ve3
wxrE05nXrrbG+iqx8UXtGdzwYBk0szpQTC4dsB8Wu2q2q/rMhTlI0SDR4I7YgVoiILF5D10zuPQ/
KsIkqaKcBbEIIkDToCDOwRVq5527MF23P4UfEJ+hc6Vopnzj3sxJvcds6L5NoQWK0zUXoskQEcef
NTtmP+yrUQIqJx0+Z6/UAlVzpTL3YMS8qG8xfYEv3/9Nj2vp9R5G13G6JEx6Sva/j+Hpxbcm2a1k
B+g78xHEZgehlr8s2jyJmFSZNDcOASVbZyi/LdRIwn1wD9deYHsPnajntetybMtE6bDok1S26JRj
XScPwbIjZynj7KnZBHLAvCynR2GQ5yd0RkXQBM3F/4g6zviI1n23wUSC2oqoRCeJr6Z79JQd+5HZ
uR2c/Vf5tF/RUAq3HJt3pUN4W4i41W3e+JJFjpXCcrMDU7xz9w7cbnTWJW5bZDKO36CLlucNcDdk
llTFMhM5ozN+gF4L997u7c7QDrcG+1bvrJ/py39IqUUA0WQt7jvOdmKDVjmIxgOHXBfnRi47HDNS
NfsFvomjkV9opQj+05XTJlXBGw9ExquDd0x6RSFlLyKLhu9+6pWr3Zj9DFFsQJBvrVoqwDxxIvf+
nvTcWDmAThEdqUFwgj/3a3p2k6J0qdPO1qVq6gbFOuEpOWjP8yLRkmLJtDztiDDYMqgrlNiSq7IZ
LYA5fBzZGsuvWPu5kxXKmpxUmgUWjRpP7QVnAxRi4i/PfDKr22KFwx+Xo1qze7eiYf2sko6EDNFG
opzu3/goHQ2abUgjMH2Gg3GoY3lODv+P9X/gwhp3i0acYDXtoMWHx4vT+C4Z9R2Tk5h5NOwkrZuk
CgT8swY3k/Xg7dKp15heaOTnpMs9AVDcqUbhOtfdGsdfM+7jqUf/8bZxz2GQe/CF8RzoCC16ktln
SavmKxU8Dm9HkUoMIA0AEJrgPQQGfxAdYl7JpVQdfTb+PazVUEAv3apr02R3g9RGl/dT9nKQgt1S
7iniyTc4G+uL+hQsPnnadc5QO0lZv7f0H5qGHGQCDAMY+Q//YMbdBJVCCPuE9WXMuKWHPii+QA/8
4mVekANdUWlVI8xbdsdgPtxo6IdpPZkM1sw8KNKgR30IgId7CPWYEgK1eMY60bUOVA4K8DRFpFxM
9f2+Ra/nlQb1IvXnEnQZwq48XEyIPy9bTlv6N6XzIKdCVQIIVnE/weAoiTkkE5qam2d5E5y4u+pi
m1oelxgQk+pLXA3MfpSFbJQo5IipCL6YXq6RrXGbB0pYrzwmbBjrxxCPUPs9R/2eW8qIMG4qorZl
0uBDmmF+QeF2HbSEnG95CpATwEyrqeHTBXTwjF9j4hhSk8eDOh/Uu7xGKcMNitFVWxopnSQ+QGk9
0Ugx6MlPV/QUWOICRU/b8bDX3LpKtQ8vttGchgDEGCypuZbliChcq95fHS3wJ7FG8xw7CepBH8mQ
ws/KhLZlLYJ0uFUIQmlL+rShZ5o+5KcGycra89t3qZUbYXKSOl7m8uiF79KwuSWcUJ1OwhJTBvMb
qaNO6dQvXCAwUXchO8y7f/BcmrBAvOTmNNhH8lApK/ik7c4Y8EqP8QL52BD4Lfxfl163g5ULZETJ
ysGyxL/FOEa9mC4Hxw6WTIzxMVCE/KBjNEMhvuq/tKqcqZeGA5CTFIuW3P4hfZcLluQzmQuLf76K
nBHzXqdEbgMrE3NLidfI9TcBxfi8nADtyZz8cVI4+12Sotapyn68cg4Bkbci/kino9KAPbRHoBaW
pkG5TjFeGIreu48aiZww3I6QtL84dsT63bK0FziH9AYIU8Dfpr6zdjxG8puwJ0dOfozjLn5bUyGF
azroJlhphEjy9NZyojC1UKezwrTC23OBL5TJjcpynKXAeyjfpVJqmuzn2LdeF/JNT6YTQhShskjS
9Rx2582IbX+z5GlU+n2isEfnZKqaHPjP/IK/jSzyik2nfPbg1eWjwojEXQgjBCQ2xFV3OGRrTtRu
pnEq+f9P44YVPtbLs3gfpitKSzHCze3c1/pfsFZF2mbwLV3PvyrnCTtl+BSV0G406dezrPBsXHEo
yLwUyqdPEWbSfi78EvvoJipMOVzxqOMHIxqdm0r9UYrFzuY1ofIRLRg7/a2B9rQ6sqXmV0wHTg6j
96izBdHq35mp0ycteUmyC1TEu05KOrf4xOS7GSM9oOPFoPTIRHGjSLRILTIlqSzoaPsLu5x0D/yq
o2lvOu9gqnQBcucU9o2i+7knU43l16nnsxwtChgL6aBb27EtilxHeq+8MVri16pkT2LOQzdjQsZv
guk+zsD2o3xM4SPv0tHFLbeCYxol7pDCP90s5YnkeiCFADlFB004j68pOUl71qLjDwR1pn+4dzKy
PIu8aiUa1dYXZ7UKbLP+KD+0xreXcd5L/VW45Slh56DJPIXQuUqERWwSZUQKDSnQQ+6BlXrta/sm
gk5jUgWsgpi/y11j2bAJU6dJVFvswmjYKMKFpYxQPHk0SV8r/7OwVtRvWfA0m5RXyREctCAU4//g
JOj6ofJ1nQY7jq07M55w8Q2Xvtx9AZIIhjh7jaVa9LQFOlti+lmOqksIyABugw9d9ChENdfmNyOg
2mdTBcs0BgLtOquh7lXJFTVkIx3hkoMMApfkINYlTtjXTJ1y+OSeJs/K9tGLxXdluDHzr3nlSVtt
UH4yEsZPq3oaBQe5EVJNcV8xIFmuG8jgDI9X9T/4XdntWMoft7jqkJ4Tvpq3H2yGyHC2Yd7Vg7zs
wcaeGMICul+7aAlm6vi0qwdN9MkE6137Y2MUacvyXY+ghbAdL1O34OdsKXr/wbGUh5iFfgRjABNK
eK4s+ci4yyv2EQQqjkpaIdeB3SBOFAoyi+4xnZvRrFwfKZU58UFmrAaTNKPOzjrXtCcxpACUO/Vy
Be5gVuDHPUr8v3LNEUQVkKH97AXWluiq0UrkvtjkMW+nc8q3rD6TAPwbrywHesqzl2UgSBbfmiPQ
Z9CY0jg7Q/0fkJZBI7x8rNuUZln2ywEcKyW31JBZx36G8Wel3C1OOJZ3xzrpmYkPrO3fNmZNbY1K
0/A5VvIC437i+CdoFtjC7I0l84dWtrbvfPkSYj0wOZnjiKfLNdnXi4DgBImqJzoMXPt1SATk2/1K
H1injynWMziCQMZeOD9WWevNmPZ23dJunPyWv0Nr1JRHrztmakQzbSKRYHYtdwwVkaSsVQdOSKZr
2epsv0jxNU961BXWFFBbzIOMkUyX8cmN+665MbMHvW72zeCFbLHyaOLkQ3XXb5e4WfTnP+2GBS9z
M3xQKXrqa0IYcBh7oIwcm0r/74xKswkr085zKn8WLfgbeV3yhBbutXW3251hVMbdMJWxV9Vydtj0
ww4P+AhWxX0LLpxNt/c4EnR0L8+8H4ddRDRvFtYg3JZ0bBS7cFA8USoy6NbmLpNxrIYJOFTmeGu4
hI+AyXQhRdiQma6By1jaXku/UU4p001Z64sln43NOrynLcUif3Y4oTaFjwcPEoYxdj0qwKnyTa04
kFgbvJKDZws9ILXSZLyCJBeJrVpo1zIn/JvWj1btr8FeVXNQEqhzhftoZX44OFJcwJg2MAVnmeLY
lFiHeU75XOns4ZyvOted/nvNV3U7kgpLXSMOsdSBLYNO9QRXmd4DM+9oDJonjO82a0s9qwNIyCmw
N/WwNADIFiwPcHBYicqtkjklg7Ip5vmI60xiHBbAVTrbKSlx+beO52GugtWIt2Br977mSo7tHqsG
dK2oU8GZiaMueyj8NPxxCAGAkzmcJEfNq/dl2j4wM7LSIWOs0y7JeD/8DcW+JFLSkyETDS63+p8J
ZcfQJlkK4DEITmRW7KIt1mxJw6yFacXq6u7Mv6inEW4SQteZJRm5o2zR1WE3xdrCsMPSYTPwZ6gu
TxcRwA/klrrW855rfSCd6MYuz3XizcSfBolIHpjJs1izh2CzjN6S8/1/mbFp8cDqvih7MUch1qZ8
AE0b/8dZ28CUQWL9oiKl/Kf7TE9vKYutEVwJuvtu9bVz/DeSVK5QQ9qiQEQ6WuQqH0GFX6rlojkA
hjIkS1hsQoAgf62UeIbfIZQSoOufFU7F5qGESGJ8w3jKYYfBR63j2gMLEWEYd+PMO3QMzqIx6NRF
foLj3j6DVYKpuiawhHEnRnw+xRPvrTifkkH/b2UvDulUscTRnsLc68uH4O+OzxElKQlh78GOlHo+
1GCS6wdqd+KqQahOeNujk+2lbGNSNflGc9XHrcIOltXb4PB8eiurVcoJ1sL35zPDMg5SeePq/j9I
fvox/UKr0joLT3Kl7VBt6GaXu+cfcq264m4mDOXi7bb9/OuIzLFRPmq8U37Ta23qI+MHEBW2pLQ+
Hcf2jkQrAW4fFY4p2jfM/xuBOWvHZEo8kG4Y49kWC4p2PS3Jec+5CjgIjSr8EldyNqsy/NYLeWcE
wI3Ud93K29OBWXLfj/jxJoeGQAAyfKLHdF3vAZRpF1RLCEikUUq2rUB+O9NgW+RF+akXTLAzI2dM
S0MCxlMyXjPbDViltpBxNT/IxB7lIUjLcQ/rgUDhWuFNO0gEZRBqQUuV+P0dhMr4Ex43ryQnftCb
pOrouqiOZvwXBz67lfduWplNkajUqMet2ABqsiaoYLTVNPnj5V/JPkeSRi6yTOtgYSwgCa6S0iMj
R5zSyVDEuRBut7EB4lD5f+01t/g0IF973Lm1mgdNw9YqyOJtSQqHDdgIFcJi9GMuApSasx7CnLq0
DGGCjeoCeoPUZobboVR5fucmlSo3NbGdYUGK0Ywenna/7FRvjaOrc+PNsyiXNTlBvifkG2jPxFUr
480OAha8S9ksUZcnn+BmA/h9JVTXU6SpVVuvKcML9sspH4rKZL7DxHfrd+RxTqVupSDaT9kyiVVL
hx6DELuGrwni2iEzUYwzPUMiDbxKMw43DqcB3V6npcLhd/g9u6RPlQ6/GHARtYn1H7Ku+JFHWOIQ
wKJIGIgPxY5uH7rakE2iJHWaUpqDY8Yc7HpVrbFjY+JO0XEUCsJ0n7DoS/egeEdrzlXGH+Aaxf6M
cZg8aTjCEh5FVSUuoRZRH/jwuZCDApgH+JXL97mxm736pUnPkmqGzgsgUNp4Pv7x6YsNZ8p9O4ei
gGqNRsAdnDH6ixCryt1yYqODul7XRtTvyn50CV+uzyp/MyCOI2om6o/1nNtNndyeb5yh47okV0dI
2jzPow23AtX87FRlpu34aSaejlqzHFQzDwwHr6c77t2jF4qu8K4Z6r1nkC3J9Rj45jtRmwWny1bY
0ifn5nxM0RqrOFsdfiKfflzIxMiS91gJTnQ9y9YQfNCeiwc/3A/kP7gWzbzIQqbKpMEmlW6QOD3A
J3Z5+bb2puRmE8laTxFocaye3fdNJruayhdPNRu212shFYvKm1+jSJ7rrRCLV6fHPXwYF4snTLg7
4RnfVGIrkqAfDJOirbeE856QtP4yjocEFkKxieuRUilwcQOPjloTLC3sXiPksnP6TzC0Mvoyb8pR
0tiMYzLBl9wtef83xvcGoalhAeO/LydUrvo719XFN4XJGyIHuiUY+fE4NmGczjd6pM4wmH37V+nO
SvsCEHn1wPBKjLsMogfdUzddZ6aoczo6NnTCF1PcTiu5k/aFogvAiAH58aSI28ZOUzVXV8rjoaK2
FfG9X1x0EJVXajFEMIZivPB4N+czkHSvs6e8K+3DExdIrTMpaIC/NWX9uzPsgpfxXQLX/MSJMr5N
JI3G5cdSDf09YNcOfvnggn7Tgb2mO+V+p7F98gMMES6bKKj+HQU1lCXJ+jMP+a+gI/Og5v+y1DxK
PjO4YAr6/ankVxzIPQ1g6BqDF46fUAWTZ7YmsmQfLm+1mdvHpOlHPP8+F11l4PZcquKbkSc3W+wk
2YqtaK4NghFwbTFkxqRYt7lNzQXNHucqzzPnZRQUdF5D2g+e07rauk/RG3YMHCmDFzufYG9m/zW6
zIskCP2lFLl3Go3+reo2wvcN5XdFcM00opY5vvs/sve2NZMO7aRn0LtAgnkIF3IZeehYmJCwvh4/
RR35uXSS9gECf6lQVQx+dGJ3x/OCNE3qQK9ZcXpZS9yEhh7NN0xMscW2nCpZIpxb4cz/WITt66ZS
rm7gr/ayhSgT6XWt7+ts/MoNUbcl7pq++33QVrm7rVgrN2L1NebhHPWXyuIn3YxQFXKrP9rGqvfB
tpsuKlXk9tn6LOfOuA1kzQraldx2v1cgt+pdH52O7YjBrsCZ0Dr+mHLaOd3woyOnjKwSjVFtpRMm
SkfDWdaQNTuwz6Zu664kFq5RRci6+LLeXDfFhYzGDWWkpDH2vdV5uZdK3BkpjFDvD1S1ChMB+vB7
v4sZxgIZUe5hOiHQ7CFxu6MATNGdwN7/4v233/HzV8LXEL53ltXGjnFRmZMMCM/f//Hhe07uuRrY
+fZZxFBXEsuVxjM2Qq7lTtDSdFl2v/n+Yd3XTR6vmsOvsNBUG88gaGVpAountPDyRXjjybslXMjz
SOVen/gAVhQ6XsEe6+zUpkF/kRQ2KRU1V+QuitLFiZ53PRK3Oa2gatayfMqHdfeAOBc2et1B3M1u
v41kChlIMJ4nBROW0UNBOsf61R+HuKu2zD51I9jZQZ/T4uAUtlIkHAnxBtPVpXiDwjk/0YV+rvGe
G1xV6RxBsAPa4xnc3I2XfAqjWHjt2Q4vjwxv2UIr+65gjdlAUppYuOigtkisYNOihesxiYofTrC0
RkI1HIfNok9NgAPqWVtQ5Z/kJ+y/D9Djtgx2hwhJ289USmf5M2EnYJa1GlZeRplajPE/Ki7FXnSH
yV4EBv7CuTXlK2Ehf0d3/P7mKVDy3Exo4ulzhj8CtYmE+G5QSN6WMjKzEPwdD/9PUyxaBVLrVupQ
M3mOnKMRDnnlJzJSNwHQomE2J7rFNYDlTFTuzfR6wRdQU2+kB6B0iDKL0A3IJsFPVWjRE93SCirm
+5NO7NLzhk14lkW90T2Y5tuLwI3wLsauOci11uXjeTcqXZcl6S5/Tz/UplnFBk/KmbTvXmOO7HUk
0bw7dg5HAz8KGquu5xgyge6jhpXESnZIDOiJw48w0LIPvXqVWrRf+RuZ5Ib2e0+qF/CRpcQnqfpd
5VnkV+ohxPdBWaLwn2xaLU2M9xQzdg6DbeQJStNrAIpOGcTtFfMPQO5qGl3kp32szEfBEtlHXTH6
6GX4UuuRKK+ZTw1FkRi6CqN2n1iU72xZZQFTpEKLa0FLfjcL1p3mEUpj7+FN50QTryJhxGD9sH99
dd/BLah7OOaee9kste8uQdBbruCeP2R4nemTxZdJLkzmNXsYQemcm2O9cOWBWIYwhGQVAWzayqap
knhWChGZtUd3of1+N1liF/iWEY2e0+cUXq8KMfc1UjMo48EqBE3NKr9Q+SD9ItbSNjLM6I+7bABi
/igLTgoLgoHJHpkovJZU+QPxfTSTNRva8BmVnENgk57YG8TFqf/rDN79U/zlCkCt/xmmBWw+BIWR
kvDK4Sf4q5ugODmzTVuHnjtXlo7+dhOrN6gj4imNyLkdoo6THWpG9CG9Hqx2rvZl/n2FMTAYvvDv
/eukvCHJbXEGC2baM4qEIIUNg4A65iABDQGRPM5UN0m7dyJJ/2Jb1AXtC6ttx2j13cEd599wZNNN
i9ou5Lb+AwNSXOyNk4R4j5av03Bw/SE4RF1e5SZy2BmBhEAXzywCmRDEv43YU0yBq0AeQEMKtqpg
j/z+jfdXOUm0VMSpqMtgAyGZGmPBfv9OkNYSo/UUfglY3pdMIHHwW+tsNKc81QNc9ob6SjtVq9pu
9uCiLwQw/e/qHn2DRxRgAU/ej6Kinseek2n7awRLTadKdAPCH5zinQ7mSw+QvL7o17aJAPAO0flx
eO6pDong852KY6S9WzCuhfLEHuAz4VEWCuWNtA+f7B6/tn3fu2Cwrk7tBd9HLKS+UMX91YhC9Gl1
nRnzbyGeeJtS0ls+GpfIpjsoA+VjpNKY9w6PtIzU7RcrtjGQV/BtNxlJQs9/ft8A83pz23uYQsUH
0CVcFA03qJv1TlXloysSo48zH5huNV8+Yd4LfGjHKvXctfnEEgk75VZyc95Eq31T3wO3xc+GoKnB
wVmsx51rAysogqTR8WxkI1CEV2K0+TC5tgtp2PHLZH1lNv0ovMiiSvbYaS5QMgdJuuLWtHtITXqe
c5iPXAmhtFIVLPIzrhJgTSxHQorHVbPMwNYz65bZqFt0VYibnJ6+cv4NG/wqj6BL3CPI1fxXLDrO
vmGDqzUwDTs5qLsqxaRHpyb1YpS4W0w9XFNMm6KvyiddF6RAt/pj+vG57w9ZtrwPojDXCOSiZHPL
DDYnaiTfswT95La+e2R4mUUD5q7bl9yuWdqNf+63TO/w+IHsvdWuDlcrR0REGmgP6Ba6zAU0+nb9
//qoD/2Tomqvf4F+8W98YgDUKQZTSk+lclAo+J3fCVilYmXP56iOPAS9CxuY6xDa9ocqnq4yFwBI
DWL2a96wz6MOrlCWXBJ1HlNTdh/d7tXUD1wAQgixNrodHwYxOOV2+wfN87a3ErlAdnMfymz3KI4l
WKbwOUT2qAAcn0d8yj1tRKjBexMy8NiLSJStJyE7KwkPJ0RueXu9tF67s/JW9w8ugMXK/M2PXdBx
R5GlBRc5ABiQ5sKw0AzLHgK7RfEWIQdbzLV2BvawEpMA2v9Aop+k3k2CQDe8KppqR1UXUyyAxSr+
LncEJJYvTMmFIBvstVQuz/YzBBXxaMoBYdv4qsc2dNpCS8cEb2nod6OZTQJF//C+UK8WtYzurYwU
K2ZVG9JjxszUM6Gwf78ktMWzn9abdqi9EZOZUigSxGevZdDizpq+ElmNiYVLOORbCNf133ccYXbP
Kw1eZ5Zx6sZbUEnuDnK/KhbAc90fz32yM8aInzPcUFbRmPZBx2geMmR4ysKAmV86eSNmELAprPQG
8fqFtaiZBQtUVSGlpEk3RCSfjFOOGXGh33ED/o7i9V70Rv5u9peGod+GmT8kN+hR7LtvJ/e+rlZ3
BVjShT0XZqz6vZ6PwOAecoCfhCAdYmgtXj7Bbl06qbiCUg9hejYc3Gj+q7I8qxmHX4a9HjRhiakP
Pa992nT6Dx46gC0ZngXBkSFN8G8Dc8kV6wDMsSBQZA0Cp9cPAj5PW5u3GkhNhnggdI8O/IA8EEnq
3Wxff4wD/ARKZvh3lwgb2EVO5cbIT6qduqS0VpO+dmHsmg3CjOAY6BY07S/adHITbAtUcCoYgiWN
0EbsGDsgfZ9TWvR8HO4xxJIP0O18eGebMpCFlHHBYHF288gk0Ikd4nOunTJd+HGFLg/OOXbON6fF
45ZW6/cThjxuc4Z3b0bxYu8C/xM0d0PabLGaIP24HM0BipDRwM/XICG1dTyhmWfbtgkfrYijSTvd
QPEn8TVobEgOd+0SGdhaPXMATNXTlTUkdlr+mJ15/xCEjbkobwP4nAOthdrTMce/60+KKCjejOqo
GVFgAFM+epCIAPNQSRCoCN5d7+88b8DTSAmUEz2JW8VCQbL8IREK+KdN5265q0mzyWkJRmrXZS6v
OVyK88mm7ZLtKr8AL29W2moE5IKyNYTDpYwzxDtRa224VcpOdQBNNLuk0lONZEV2pYbuO97cC5cN
zardWN79RVY/f+LDPF5h6eAt71sFWowO1rbnaLGPdm8+JydH/0VG8ckreTfvphcq288hVAAYTJKH
6XTE3qnqhHfP/HuQJSZ5z43fu//jatgDjS23XZm23ZSqBajsRJ9T/XwUfjyjUq+P2I+riFXzroQ4
BkKzT7IwgPBdf8o/ZMciFdZ2fAkZOPO1lTNZzjMErRDuUPWeaHx80pLbGRnxXUp3orhGgenamd66
qfTNbGx7KdIoz6jOOCc8rmK4p6Ko/hKoACPagWrXPg9w5Ncsfbp+/p/Sl8t8ZZQXewgT/S5xmH6u
Oom1Br2ZCKFVaedqAhIOKlCOqlUbfvXl24eATPB43AwSnNAGd4oAE3HnU/8DfO957Gpyq4xzodvz
M54Us1nh2FVImoAPuIgp4j47yzgTr42kJaW8xEyzqYs7PiqM18tF1ynRpRbSiengc4+RCFIvGl/c
Nno/zY4Ak3U2VkNszO3BREVKlHuPqljGwPm+wN37vyzx2LAzkfN0EWrJAHKiNkcUInHf1cs8pBT8
mNAhLhRAy7mkS9TeSRhR/woT3pTeU45Bq8+J24YGJDLVywpJB1nAyyqf41gZaRkjd6GIe2nixbOi
78fbSy+wFW+/kOZBDxESzhu5SdOsiFUXeoJZKy7YnBsbYicYpnY6J4C/PXDmzjIFdK7BOBv3Dr6V
fxjvg8/IE2DDRU+2acSvZ+NoZ8fWz4TH7cwA7rDsup9E2e29/iSEzYJsQ5AZqhbZeoVwSYNFuulu
RYejKMOgxSNMEjL0ARSjclo6vsGgIRBLorqKjLIVjZEypzb9iqGagwBll6zdJyUSWgZhN9OCgxbY
bVQPdC+uOLp0aCFPBvaENDepO5YWawZ/8fTNT02XHx5LQWDw7n6I/vZmhH8jdMLbJx57eR1X0dsi
n9KYHzhVYo40jYL1DFAxvOCplMdEF51Q1aHKjVnXKHMP4C2Mq9kv+LKHmAKFrXzYpQUVrdcT9Tjh
9db+g8Jh/qXgyxrXzy0tlcknSyjWrX6y6V2dYPvASjAXKmeHoEkNfuqf5dY6ZJcGjRsgdRSerzIB
FsBllq0tSCOceWnts6qhaZ7hSmsnPMFzqMcOXTDPHBhTofq41ROucBNTaOfZ79QTmWmImK2ctTns
sxsYaSZuvT+p3o7enJhgfenUA5jz79rMBeZk8sm2Osvf6XqN8JeXpuItG+xSoeTLEbPF5DCjjH3r
0qli3ivGk5LHhkt+nFaRld7cl7IZpQiFEvIHNZX5JS2ak6szLhjdFI2uyFAxVeZRmpxkiy7YXPYe
oYhbHyjdtJfg9m1O2aL6oaRVrIlpLNTg5q/gIAKkvI8R1wz4SueomBnOz+TYwH+2Qxf8b5tgQBly
QWmB0jTFXYxs0FCtXkqv/IBvLFwxIV0lAfZTzRLD9IKOis9Aw8DeGre67Ekeqp+Wm2FaAnuxzCAz
lJzeVqXmbKDOy2dL2tR0TLvGXQjM2dIChWlZ6THThIWu1Dt3wMZQdk2Q4mYl7y5j9lXec12pj01s
3iaP69ipgcoXQrtHOViSlGIysypKH+0DMR2C9Kp4GyeqaQPN0aJnQEUQeuc+MvTJXpJKev9FguX3
XTovBBk8XAGf5QVvlF6tUyHC//9J+/1dqqr7ICOsuakdXsG2TcYOSWd+FvJ8xMVYr30krfIl43Q6
KJ6TpUqAiz1GYZcOSHdoLmDGsOMhBPK2b3yOFAm7e24TXhgPS+q0Ar1QBL/R1Ynz2kScrGEjZwCw
TiIH8bD2O8Flr6eIGPd7d+uC083lFOgSzSf2XfFuhJdOP1e5LpOwOV9PGwWpUVcGIghRfJCo07VL
yWcUOZ7JynPaJ1z8Ma0d/QqdMAGwUuYBMQx132K6KEjKcv36L4MT8O47NgrySdLYltZ1bHMKa1TC
ljbd8uc/HAWMvLo6qCT/WhAbjb+lysfVcO6KQKk5lHpJnyY7p9MR8AuxI8o6wnWHLbX2fPnwyO3u
6OjfZfGSanxsIfQ/s6n/eXZ0OGYC0ZoQYnRhPHnkhKjtnCP2d7iNtujyZ9ztjnPNl5/X0nKOzmCm
75/3fSai5wE1D7mL89AE9j+KAcK7YTb+S48ur3WbIaKcbUR523t/7iVv78uCwQPQIMbXfVCW6qFH
Zw/Zyumy2Lj5d7FRGQyw9uUwLnTH3JYQUaX2Xi43iG0Ue0wP525l/NklTayhlpxhM49u2qxVGY8w
G36ud7JBKowALQKLNF9jaZ28SidSfetOuYyDH7x71AQzMLIwuSmzgOVzn/nCsLJi3WQM0GyM8uTf
ZcedaZjAjVv75MXXVuaXBhEnvv9bgbQqYt165fRyChUu1QIZbnpk7sVUdsxZmykPyLFIm41a7qrA
3/xGzUUliAmaxMbLnX1D9GxDxxxBem3oS/UXS5rFwr6Wo8a/tezoOX50v8MpbeJKaP8MnkFLKrs9
roKka/APA2lCmAeQS5uCpQsk1ZMRRpufUrke41BGjzAyPTFvKmliDnVlNC9S+C2v2jjm2rzC3blU
UqKh2CSVsQolgXr69Hrq9p8wXsj31gWJepwMoXW8PjNs2d6nPwJxNYF+CEUCgzRb+oFWeleVduOf
9U3TT1WmovRfLQ0S0Hxe+sIxZWjpTkuvS/4lJUFgNZSt0yznSt71UhBkdCd3Bm8ew0j560FCfSQM
gZfT087e9KFiD2b8252nouZKEVOYFjbha+EzwcycY/vOTLRTSvlDBka9UnCAeICAyfp4Qz9mGGPX
oHO2M1HaWJMXuIECdJ/hBtmjsTCHF5lGz0SXjtEbnxuD/j6HHpcoXgcMejlGdgj5anF7M7KmTRtF
oXhQXvpgxPU+DHDqTJOwTLijIp7I3Uv+/+QnbWlCfJSpSTNe0Lh9iiUCFINprrAEiXX9DZ2q+LnI
iuiOKfY1Jf6rIG2IrYJpQtaj5PqkYaYmJjYUG0tWjb2snV7AW+QWQ0YaqTf3ApZ8PxKOpUSpjk58
Krfus/ll87EOfrVVw9ccSxu9Bwlf62lt3hQnojiKwJKWQcIwDt113GmN68ptOIqX6SSl6dqhlOxi
E2iN2oUyqFExQMjXD8IPL+5hNrUisCnDipONSv9LyWZ6AAaki67bftbdwvHcG1xsCKAYpKBSoKe7
PVwvH7nIgtL4atSwJCg5OkVPQyHAvEhwK0dv0+VmjrCPSHWJ1P+LcZmx4JD4XL6CjRO3PQ37HTUq
y8C/+d0NchsQOd3Fy5p4paLsMnflG49FNugti5NRzlHVgWvSTRvxfs/MhSvzGfR4m1X2ecHPeoUZ
IKTul6tZMVUl/L+/Mtg5w4+PPlXa1ocDHK7U9++GWebvpT4aFQ/a41OSkY+CWdQyN7SQ9h08xd/X
mO/oaw5gzHzEQoD2rjFL56I1o++vg0cRV7SVeJzDZ+yB6agFrI+6Os/4uBeUj1ZroRE/qt3b0tnG
sOwXRMKfZBiZAaZ+otZzYc+VOEy2KuAqF1hjfZG+CCr1UdG1hHNSDx+hpiBOmT4WwuDkSkjkPIw4
UUDTjvhy3hCYFNdz9SSMFIaAdxY9tTnofLmsEyyNjnIrjvlhG/0NUf7A5vPjusRUpUvKQQPVFZhx
lzP1ZEfoU344DQxDn5fpafgLwu4tVU9jFhBSyv1h74JfXvKFRcPSg+gOXRJcpOGkRsBJi5L9kgeN
VoykdOwEs6nC5Fpq/VUTqgKfHNWvRiw2COhajngA+fTPfkyfKfeHxH9LU8+dE26eFrOzJiWBlr4o
ppF3eA7gC+Zj7pi0ZaSn6SaUodgxeiJv/Yn2lALtVHuhA3tluBYjbxvuAxWwib6NFwYLRbXHhlgA
W7LgybYFps/uYPcUQoeUXfUqpjIhIdRSEgEvE9Mo01mOG4EFKCn0WYIUqexunF1uvzDmEwlDw2UA
ZA9zKX4Mnz1VZxJ7VSgK4ECVq+xWRbywArPdfwps0X9hM1KX5AohK+t6fghVdTsGE710fE6+ik/c
FgP33EfoMbDcyiMsvyg9GhrpTil2punjqxwnZpBW5rhOUHHXjVL6QVSERI33oc30yIOF4HRcpv4q
xxF9zkeauSJ1Hu4Wyjzt7DAlN4LqrfkPHxu7jajgOBdFLdkbTbw0NKDG/hS3oZllF1m0hTk9P+ge
weEtbz9mvB12JgvoAlWkzx+qWjwshlpZ6/8Muy/XTOjUZR5dfzPaH6axAc4hnh4Brj+DOst1aQpR
zaDlSIPs1gaHFohrHUER1WspBCTUuQaprkiXvAI1FX8R989vBobgwZPgGDYUth/MuwEsB00XvohI
XLA3FpcMc0BEZfgGCZA2doem+oxUIzaVp8r7rs+Y8gT0/JOFp0bzandwvuNPz19c6TN+vl4lnEwq
XJR+Rg5jZRIH1Bryou7Ee1tukf+FYGFZREcR/wpFFceKBTcJ/6yd7kcuIEO+F2gKFo3vrFZeXmrj
IKDrz0G2AAZjXz9kBgwsSYWME8/LLdMrKHnvR36An+IEfYhIbCDZl1FHKjHW9lbijsvtEvcVQr3X
t137iwD4vg1o3XrPmMoi0q0ak1mXFYFAeZ+L4GL1ERmvIF2dQysoCQ+B8zXlJk2apygWmu1y0Zs6
KCh05/uHDzQUKznPwPzBwO+T3ZggkEWIbf6OpezHpa58sqYFNhjF7iJe3O6KeyGPgEH3WUcczMir
oZywXQoMjzuLCUEPL3QsHfDuIKYm89dwGnUg/x1Swd6h5zqMa/3v7Z22BqryP8bK9a9V/SmL4Pkz
iqh2VR3CEYM44Io6ZQ3X/7cdM7orj5cTYcnN96Q0DjxTV8x/X5JjJ030xZShPxk+V4p5puIsL8Ot
pcRg43IL9Dt+GRXkUlOjLGONKsZQjC3oj9dVmk5QujEfrmjkoKdoE/ZeSBf5vbPNO7if5OHSddAq
wk4Bm9FMxrhXkZsmLNRMmWIssG4/tvZpdILeMtApFnqBh93PPBtVJcmas5+87P3gnrdmXAwg3FNy
WSE6TznRpNtBQGxWPDCDkGSl3gHLl8H3NbSdzK28G3rFG0yoPEAEwLVjXFPB41ALtqr5GkV6jvho
4VSQ8F7luE+oVyHtie7mEDX5v3ciEfQF1fO9Sx/cPdxPO8y2oFUvevAZX0nqMEt1TDBOsmE4DtLM
ewpLYj0csWrinuBDcgS7G0Hg6i/GwnlYXuzXMRd+qHgA+SwOi0vPpeivaXBkUsOhSQOcSRE5OfIK
ujnMNsO5II0AC7Sv5LvLKqrS3E+AHgaEeJdKgI7CB6jeA69VA/V19FIbkCp9xjGsJSa/v7exdHsY
zu7O/N7gR32dqzs2EvRBBvJC/ZTJFl6Uc+RarMdzqmk3KIxVqFv5Gggn8zcN6PKQeWfxK2uTLNv0
GQcTZTFUalJGOXEnfNWXXlkkQxfdUDdMjuMy4BylD/ialiN40kOLnWk/7ZZE0cfM+8EWg2N1UXv6
NnBo4H0Sv226Ry0wKxidr7s/n/Reqq1ZoLSR0aHD6G52mALGJENRTFDV/h5+ConlCpUXHYDWxn/M
fMVcd0ew+NviY4DrBWc+hwluZeZVzD/P6x9+iGmFBjH0INaYRc9tI+bQ+awV1wad8z8+ZwkSHxBQ
rUdR37Cxt2d56rJd5OyNkXW+oJn7SzBoHPNX2BSjBabmtuz6PlO9rEHMoiwR+FkNS6SNO0kr0FWt
7g6OQTurZVWRsp8E/rcJUe1Pv2dPQgADBasmMFKg+6EJoplLHwUDwMpwWEYYfURoLvrYeZq5nr6V
iN7W+Kitmx1IMudCYjLjnSs3jKGFW3kL4iMpHKZq0REsRS0F33wIjyjkVtpFyG7IZ/X3f71MPyJg
4y/z1wx4ef3ODPK4u8tXUar/1YfWgS+seLvrZcosX9l/Dq1gqUu2/zJitgVjKW8ZkkKW4cGFFdP/
2W5dwOk02Q7ctkv/OtPpnHZdVuRxzCYECPuQ1Z6nPve10ZXUV7BdIJaEs+QbUA2+gwN96tMNFaq9
b3GqfcbGkY9yGO13PsQ6zLw7vcIUQVs2Ft031CAvLdoUTd90yxcm3zyyF5B+cuNssM7S+elhByUG
TLVkpxoh3ohHoh3opRvNWS7Vsjppj+s/akk+8sWayfFb1BTRm6h0dwaQCoQNK2gUzi6m3dR4O8+V
5CeVuIPdBnsBeeX+EXcufR9u25/rXX5rNDUMNs0Ljn/tL8Fwc5xrPj4uVJD7VQXWI9Jc0pAgSGPc
Yjw5WxVH4OpBRqY0hlhzT7n9N0yb1TpTMmQ4TGd9L3vn/daNXFoN6L3V7xwKALJ9ajjq3V+uEQ+m
87CplaDD50t4qZh7YXhNsXRQXS1eOv2mj8NxM1RjD2jaM2DU1Fb3qXspwr6pfzp6u3E+0MpQg+5K
IKRDEY+B4GVwwUh/OH5E8+uh//6p6LbZ6nUQNWciU7Id0ldNS7nijEdnmWV8hFrzJOLRDQk8MAsa
Fu3RwIKiJ7KMml8KsnpL0hltyXwql1xVXhFkTQIS6SFxymu2bNXYybm7GkG5iFywo0oFLgOWzWgp
5M63Ah78t0AYn61XIk/zmCoxUK5FmOi47fyNBiNKC2+Dd2m6v+Jxv3drtEEKsKU3E/otzQPar+Iz
WwqvwsYzuh08zplZjBRzrng6qLXi7Pj6y4S2dqYphIyTbiMzudRHdlfwGgXysfTw72M6LeLFQmxf
LIVa+xOcNnxHm3bEPQXLGXO9qi0OkVjMrLtAqPJXOWmVaCr6WCjvKCluJ/d0RLtu8TnU3Uz4aPoF
ivZhGh7PMvl0Sq/11bECs0GcCO8NoTK+VzE77oCpLLZsApJZeiyUVshrvTitujww4ACdtUEwLGC6
Gi5utkIVqGD+YjjrSPAPVl+rcUGenueJ+KMxNXWmOn1SnadgVd+J6+lmUvhNVGOatnd84szGlvfe
qiqebzh4VRA5ajDpI2lAcCE6mS4XYNI2zuexkSiNNzTDm8HihrmZ/Pk3Llwb0kvg1Hhaj5Za8V2D
9mXGoadOAW8kRgH8V2/lUa2N25pb0RG0HS6GgCOBHg/ls+ubMQIjirzP85/vfQOwNw0q+j4hYg5W
2/T19JWIn9iZZZveWrvnXBLTsXck+4TBBakdmfh4jNDEcaByppLJGDbaJSzjlLDejylEkDLcENtQ
Iz45DZ5Q9PoumwWZdDr7NsGZslY14T8JmLy3HgsJpD7iRLm43aYYuX+zLPNrzaRFRowMnJEKAYO6
VBYqfMarZ7yXwpesA+V9UTfSyLp4KfXlLQpFZKuNt74Exk8W+1bRdOhDqFIaKNoVZPtckYMwffo1
57LFvHlXOfsaKWAYnAhYzJoaGs+3XYEM+0OSr8aKqjUhQAlTOsfD+34eW4ap+xa5b8LnflKSCdqy
rd2Zq2lUpRdOFCO9wGP+WEma/4PNd7FzzNMIVnUTKXgtEVuay1b22nC+MKWiC48c+wyx8ORSQhlM
XEsc7IGZriAuAcJ58C2HzXznZ4PCbqO3ctYxmtTE028yT1VjWAa6Oxb9gBTa2v8FgP7Owrzf7t/k
IzpNxGC20qEEIGwTftR9xffTN83NPgp4TDgXCETQjLZuXKn5i7TfS1TvpxpvWf94nHvGyAVEsr5X
bXAcLZCDcDwF+4zZVHY0wihS7rej6/f64PiQL1CNEfd3s7TB0D5a9vFXf1ba0+4F3xJhSIUs9/dg
7y0QrM6f1fe5m0PX6N2Boul2vMI70mlOhVbzSxpNwsTJYNioXWM8U1TKwAqi5VmDTX4kuD7YGdyD
n0q9xpUT/1VS1oiZH5yShywc3UggMCw4/2dRV+Nti4ze8kzWTLDVekNMNd4gW66569uRSmLvUUDV
Ksp1URfgF31B6JmUHCTijIlpf4pps1ospn4ioejwF0GdIacusbqODeLHTNkGzN4pxOvgXSGrNI53
fiZ40gmnNYCd21D/j+OTCqQKA6l6N1GR2wQS0fAZ+w+84aUtXHhSOBNphh7pleHB/69czsZdhtRj
gyajS9K9qH12xWvePG1aGM0MEYM3Ea9nAUQ/ThqLD9ipdj5501NW9sBBxpH3myMf3RsreY6LAEI2
KcjVV1e0LUQuSSnLHhfX/S6uJL1JMA+pNBAzp4hWypvObp35cgnSIjeBwZTb1NKimv1z9QgkDexh
4WhsDW0U0pMJcMJJG/QdnNB+/5fH9+XPLgaW1Vpanfj1mHVoYsRpJ2slbKN1e0fNfht1TTrdMbGN
zawy5KqiSi4BeEe1L4DNW/fA4MsFR6yPZd2Ss/sy5GK12rUyTDPQjGhXaMM0AG9IM0OSOR61ZKyo
rG9JaQWWRO3Paclf1vNivRQpLjDR4ezYYPbQ4pqtm1/IuMLeoZUXgb1ny5Vsk1gURr8sKfsYpWyj
/URpsoo2A8u3d+iOpND3XKnJpzjVYRpZquRDsTGxsabT/knEN5JT6l16OOReN6HOK3Wi3v+w5my2
0ldlkwqJ128a0KLm8JWTxK0xPuJTku2s31Lr3mPewYGGlkOK+fWuGP4e5hDvOoFuk8tCkiYAeA+/
T09RXR/G8j+LyFOYU6bYJtkyk70qXiu7TVePAtvyz00nutCDwviEmmKKvp0boU4SIBkstXRHZBl3
p4RdVblWEKRuCrNFeNBPihday1HBdf6nGUnHFq29beL9JYZCrqIqsDpHOaRmAs1zyVbVcAUCuvUk
ndvj0sl67NWfMzukEHT8LTF2ra934+soxs/FFHpRarC0gw1TSU37GS0gmswcAp7Ocat4IRHR9aBb
PJ7OBzunQUbTYLWptPuzim6WlbwHLsyR0yGDiimumIt88Y6IluhtUNpD+MRR1QcKMaX2e5URXOgz
kEDhwBZHAngE+6EZRFJ3n5ftxg41VOdkRBwgtnuUldApWN9WIvgBzJpmAfKXtPGGcwpu/K6WudbB
wf9XNzd3ddtGTBGBg3PHfIbFxLK36rR8qIhd81tjWcX5+ApwytCJ23RcIoEwxcLEIzg/3OjQZd+A
zF4pPsMV8+lN2wHHPT+wRTaRgV7oqn1HLvbe3OxjyNg8jhRSBlL5/ZnGnIag6pyb+eSeLMRuh9qn
8HsT+1/2fOeNVamSib6fJzsvXats+oKoRkmD8zYKIh1TZmCAOTXGRg9nyT3xw9vlHv2Tm4Bybxf6
g50J2ZQbbs3muQhjMALZyffwBDPwSWre69VeQDRFIESfHab8pZM9CCykhO97XbP1mYes7hpSR6rQ
abGqU4jgwz80HVeEd7D5AnaeVbiCLullw+Ar7lo54GVwRuKSTY7M9zo03xeDCNeqBKEuZZDN77yT
+Lb0gXdViRXKVQX/MupusZP9jW7RrRzQXsrovtA60V7VRe0nF0djGVsAVGeGohjBCJT8/WMqxEDz
Wyiky3xlTQ/RjR63IF3WnfToN/Jx0NSIZasRiq4Y+/qLHis/rLWYkyRpg1P1lNTQi3+gKGPyx27P
PQquGGPSQBXmP067ZF/FkYo590pU5Zc36MAwwMIz4j4+IXe/ltBe5se/PFgNCufAghRZtma48rpg
Da95MfUM9zeaTiOXaN+5tNSjCYDut3I8d+pFcEIKivSmHncB+sO7LXMmPHagJeY74bXu2V0QbpJ+
H9HHFxPNkQcIRV2fuVHZ6F5io0SwtGhDIiTE94iKwg91QTEAZJFTt1VDfZ+N8o4hpbXQnO8y5LU6
ZYnh/HimKxy7enQlkPL1C+kkvX1+P/gWcPq8N7HOlzNuRvPAqNtADOUsRbPNO2ebwaFK6+j8GHNR
FaOQgPDqMUqnHMdchiT2FOksvJy7PG7HlFYUDB4/hbiOPGXMZUFZeZt51goJRVtUNmBdUpfyaX7W
Wh9xKXIgDKrtXcJ3civ62/XGfa9JmnpFb1LnaYrTh6qUglHOlryZARMVlnPkFQJoAsGZ9SHRNQwm
piZDUl/lhnKy43Q/Vd73r88pzZ5dCl6KXZUeUAsLsRM7DDMuyR3TIQaIeMmvnRFoG8Ii6uGcQxWm
LtLFYVdcWZnkpwz88rOAaWugmdzyHsRBOJLd+H6uCrVMs5W5GrLhIIM78iw3vnq07je7wX2L3jNg
3yYDMyAuSHERVnum6fIV3JyG6Bvo/2mNP4Q5ViegMa70UNGGtTca9hNnRXbGSJpoexqfc3q6aSOt
NF6CbZuVMPA1XlqO0Hu0gWnFptxcbdrEB8iz1lzq4bubErCYvN6AkRWTUC8fHUM5WqQPX1LGWCb5
grD9cgxDEkdHFIX9X2fWH/h7WpQLIAC7gFit/4f76LAsvMDV1UWPQ2v1Aht0Us8Af0Xr/vfZeUor
M4qrDscTn5WqBDlPWT8VoW94N0A5E2dPqyWGP1tmSA8tMl7H6wTmC7AwOAt6kdXTmrFm8l/EkwMH
rewBx4Wmh5dt8BRrXRvCa3nIgIlp54VUU+qF/0J7tqnypYx4oqJZWxbwNkZipMwU+MH8ugfOHBmd
M5E5e3mjG4nw/JnI+8w4+cRRo8R+1HFz0fVw6JbygcqOJa20PA4LYesOV8qnhSk3iBsihqocvPHv
9UwYBGeNoRIxNgKAeZyrrXQWKkfGAP4Zg9F5p7IAhKpGTSi+dkvwwukETqU4gQH8UrJt9zMveBbk
Lr1AtVUBCNkuLJr5azn4UaeW/JYAxFN73fkqhucMb9Dzs0l9HChLrcXqs48gH5y+1t/5yjFknVzx
iTyfo4rkoLpJz0S7Q57q166Ii9hGXRfmaYL7i0a6Fs6dtIypW18V/1gZK6g3yduJWjqsD4s+3l6D
l+bBr17ETJpPJEMIPY9t19oaCloPYUXji/0xV07pb1n0ulS64dAn3756KbJRRIG7TBS3ofVinWp6
18E5RZgmhTgdY0nh66Y/4tx4U/CQbgxjbTW/SCoBjfBFkJ1TFxBJGoaD3iriDwLOzbLNmZq5tZBJ
XeRMUg24fL7nUx0vnSa+JGdGbObaUYgnh8oz3/LYDuy7G+0wr9BlUlUawLCut4D8pHX56PFWGykF
wJZLKZykG6TyUtv2ZtA0xx2wQRrJkl+NNmX7BxWp9VimdRsRlYpNsBjsdHTp6GELA7jEirpkX3YX
gP94G0MXaDEZStUFY/fUen2LtIn4JGfB4obS07lDXmoj/vL3tOu6HcKuznu9+6W7IDs2OLNee8UP
YGZuWcG2xMacF0V69Mfr5WYvOytV2ThUk2EExktcrQxrGsmGmtMWECrDOd9slqUM0BbKz7QWXp3x
4yz3rs+MZsdtTpbaP5HxcrqSLSBthynO8IeV35nqj3NpCXera8VcwAqUajeCc5NJ1/Zu/z5T+4ZQ
p5USZfshNyY7U6xmNCTG1eTP1XoPpIgdEp0lt6wmpo4fe74ymc7DlMaJEvGsWusC0t9kWcwPPJ5R
b2NInPS45l9KAAxSbrouj/KXhgbZ61/hk16iybO2BhH1E8PBlpC+e+Ew2v6qksLZQV/c7VY8N4CR
UOycUFNsgsPjpsQNosXMr7LWgPNRXZgx2T5u9PZW6pygqNSzZIWMKDxTy964gN28ZukqXBi3NmZU
BubQHCKIWYyJZ4RUJr+R4Cv+403TFqOjNly4l9XYyQ5zuGEl4AsIbhEEsgYKJWfi54m8v31v8tSX
LcXXyuov0Ta1j19Xw9PlAMQVUQ9TM7EhhRg+yzFnVjd1IeE2atrfq2auHP7zxwpF5Cv3iweZznUe
wWhxPGnj/2ibzKUxKlarSwR8mtOAau99xnbgSDZspHsuNV33LxH52kFROE0J6ViTuQhDtzBHdJNc
AupFVFqns0f2nKvYhwpF8fXJCiEjIEmgoCbmf94yFIeN7RyvMem0lvpvUCxf2258vuQIcqXU+cRS
4SujP0fKHoiks80+A2DG0QR1narT9gtCd84Zl4NfYvJOsM8UGGWdk1L1XZxxB9u3QAwIjj2zZpch
D8aoRZosHTHMopOWn++0NccRNKs7jUfQ4oTWJbFd12cBEA6LQAJr326cQysyd+AxOU0k/6vIVVbn
nV0WuBPTWgFDLtnEGsNgjzlmJU6YQ+wvqxQz3VgJtltK46x6uhCuwCmiUurt+U3bwkk5GtRx0eZQ
MOk0W+CnFY9Wlvsa8utriqbQswrilKx9T44nR00GwyXms+r7MVihykBDgLtiHMtxjEhO8nTBdu0D
rjvjpFz4t16KI4s88b84iIqJMjxfVrysN1gkk8VtN+XVTwXcG2MvWs/QGihGWTn2GysS6wGJQciG
vV37ug7OagZwEYj3/xLlGg5RvB4bb+H/2p7FHaMmUu4+cwWALC/E69nlRwanrNzN9jacIxdTpUQA
nEwq5o9eOeZqYiHADvBbkq9PIBy54Zn/2jde30o4qqBiBpn59winP/KOVh+Nn1I/Bdkt8K5AwJP1
aNczTU1AdJFfLN03CCuiZRyaOvoCDW2FezuxGeB3OCE6vovo0DhQeaWoFAk0NP6AW1ynlUaNw/yq
zBrhgspvaGtyrktz3rhtuLbj7+0ulmB2j9gzsS8vTvnpd/I6pkvvjKHJS9yPq+jb7QDsEYD93+EW
/bbjuyJyy+K+CMFuapsq+qkjMg8q6kANV0VRX0BpF/LwoN38L9VFGbxC2Jf/NN+mKkhQBxGXvrWH
hOtBEtr0ea+OXsZ1AqglO26mUS1tZrmH/a99FOkJO51fNgRdbYToP7uszkhHrk5LwhhOjnLFvcTV
tj/TcpD1RCaUbR0BaokrAZqnNy+tLYvrSOjLgsKGDeyynkbqzeB0lyly2sJgSiobyK5h5Ss8Xzdz
x8+Zp0LxfsrSZ7KcJ8K/5qzTLu+b+fqUuHJe+xR9ArfPdqiBb+PS/qOdBbCaHVvWCE83AWuS3GA3
Zs2e21/PJnA13l2V1iiHFwxVkS9Rb6RRCCzP4F7nVUyQpaR0CJxNBnSoag2opehrUOnttNxdn61K
KxlbxAy4EP+qPTEglcs4JYXW87/f2VhDV6KuRCGgGnTWQYFqmLOMcGEYpRSjZziCSMeR5hFImZDN
1yDdFLYTkyxtmUlAD9CJoEeTV5eTAaWPBn5tI8e+THbtnweRsxlZp9tLUKwhpvpkUZSrp4m0i1fj
xtCQeHi2Sv40johFppjipSccRbH0zvAwvk0GF4rqEziEzcT4MZkG9cRdRK0WxCU03RGMlmgXxSvH
9qicL1ihsyCgES3yB1ZNTP0z91o+dPsrQdFYfFa64wHOt+4b/T/EXW2gPSuXVliXy9Iv00l7FUCF
N6wcLSYEzA1xJLzQ+0Qyi8EY2vnSQN0M0+tJay0k6MSVDw5e7G0xcUx5u2/05Zv22+j9znGrR0Jk
Ororgr2M5mFIWyuMSbXcuQEbuRx3t7cl8/eT8+b4rH9m9en8NhQQiTqsuqToCxynJmsMqqkhTGZZ
gW/N+g1/NvfxruriNGJdPn1OztqXTCS0Sm5QSswD62ce6KL4l0YB3MtqDrwBPaIzzVHI62zS+RWz
kPKt+wFkKy2sxNwslsaBD0Fyj1/yv8vXgyX6pXpjO30esbKlIhtTqrhGNXzweHgKTv8Rkrv3d270
4eezDgiTbX4ri5Fq7skIMO+cszsgD6VkEULJkil6QI93ejV7F6uGVRyYG2l6m8IhZj4nx2EWPVFE
T2BotO72LP51MqCtoB72qp98rsWWPYbh+KMXghnoQ6ABxTfZoXqbghTIC18QwWxpUxNsPWxihNtM
IdvPCoUYkJNFO9zVeoQUOWbvNioseKhdmzi/V17RF8NGI6gz79BbBWptgiJ2cqYg+C8hZahPuPXo
ikMQj5j12SSdTDYZ9IMzJ+OVwpEIMtjVuMCU5tcBq0MU808MyHtayzsFhIZJoIExFBfWtjceQEuy
2Z4bk20kIblW/2Nh8SF2V8t9Zt/FHhrOPJYxI10KjFZC3f/MK3Whq96cPeqt9shKdFUs3bxK8NAQ
bH3hGAprhfmrh5Ffb2xjkBH23QIfkvHF8NMnUnReHkCZ+JT6LR7MzYdPKRjT9FkMTl0NIun26UMM
Ux6SmP/BT8E38XvyhtkzzGOhiUXj94uSMjss40nFzdYOCTwxKHOOp85RTew/n1ijVfzoS2F01Ckp
FrYwleb77OqfzEPQ/suDYEQ52oZIIvGMj7iyNLzeea7Aeddqc8J6wtE8SSoBsKSSfoYic+86Q4PY
CDiGL3+j7LqSjF56GpGM7bhF6ZW2IUIIxX5rUmhLwEu9z0yFIZqIsUEBDOAhtcVpv2hLcVbt9S4J
EIA03s7/SK7NqAf/W9br2+1N/NqxuzXNa4hos9yjqlye3I24QDrGigW6I5N7FuVxRayd3c0T3Ui+
63iawmF5wXJW8VSNcMOxGkWr8yt8e1HygzJKRLzZhGQiDdNBdbogCC+pk1z+GI0L2S3pFl/t5jOa
RZCfHxM6a1AcyZOEehKV3t97pIynxE4Xrm7wP7yR+QvZGm87PdlMlAUWhwffIbI3qgU9n5z6JH5J
R7ivVgk3Ng+OoTJ3JZxb+eruxlJNVI8hkLhVl65WbTdqUqj0y3xnjwfe8SBH/iUA3j9VAQ+DOgF6
uqDrq/qwJPEQJ9ojdEWG+xvMpWc2y9t1gOqTV8sfMvIUwRTQQ/YMl+ACw6xgejmRl8Rxm02m/IBY
XTUOOwxT8pyFN+A6gt/okUff0Bnibz/GIr/9/GJ88ZM/wpG1DCYm3AtfRauomIhNfzPIMTAn6qUd
lEmU+uCImH05gQwVj1ACLbtRXtLu6pXSdOeVlNTXW5XaNGwOxlzQzdpqM7ljnu1xtoTKAdyr30t1
5vz2HE31DYM385LRXeXHr2R9BOjc6a2DKN+pS9vcyABHpiPJk2Hbx4h+w6jlLnwHDeCaQAA0pP/U
htrz0tQYgWtjWFpTd1/bgs3paKYotk9/qevrOJcwSxwe5ZFsZuMBzQWNb7UAsbnJjFJFgOlwQ4ti
X6Llh2UcZWemxI1eG2JEsOLHHaaO5/nXjWjw8ZD3VMcZmctfTYeMBAqlDtdXHm+HsYTmyM3gLHVn
ncRfiV7pKowaSoR/Gsu3tuXNyh343Yvfr0zA7oK45vweYuYO7SvK2WL4uo/IKIu+ZuwvySU+djDt
ryvQzPpW6AE3EHqRXiTt1bJ1X8vcWAhOW79aHOHpBRTpZZG/Cy1U5X2mAKd85QmriDQUT3v+FsqZ
2PLfGT/d8dl4VYVEI4XewlGuRoCp+tDPsZ3XUbMyhSP7KcJHzwusLqLIEDap8lRM/HbScrNnfrNa
LnmyuK1m8xSzL8Sf5rcsVBc6vc/wZdOPEZHuBFj1jEgC4SxdVI8ufiysBRD3iw6RQODtDSbawynx
7iBChooPWlTlPpENm4gOu1D21rEbGPuL+QFhRLkUM57EAwEWWi6CitZb2VTq6divtfXg9yuNVaIf
09/H1HG9tlEBKKdPdyJxGe1QbUisMA6ObzfO65SxHhu9UHmL1v2SOrE3nx+6/kWiV8PvJzMYL2xr
PZVssKony1phsdk3QJC59EnvJW/tMEsEkK4kKJ/wh3sUfXxKtALLi8gpoalzxiAA/4OsOKNQXeSd
8YgJ35rK+K6e9jcfbWlbc4mRXnG2ip238786HNt0FZUhboY5iIuMEfk5mmE8jqfIT1fYmxmWW9TI
6qL9DLgphRYJHoGlqEAvDPl6YEdeWFM1pC38YUiz+OyzYkBEVmHMrvI1xKJNNIuGPBOMpUt/A4gI
M8zblyJSZ0llHM+a7h6zcjoXUBtgROB/67ysVBHb+EEruzw3LHh9Xq79jYMRkDn988skndKeqkwi
0F8gvJNJ7Qhr/eEubhH/VOSdnIiyuAjwCQMmTFNMs8KVLmpXUIfTSlMOtBZQwcx94I65a9HEi3kC
oyT30YijVTfT7rg0gBXgHRf1WtBSg8fx5f8Tx3wumAeBzH/IuRjRGW4OGGWPF6x9oY93J9SEXpyK
uRQEWK8h4QwyWE06Cxwr9HcHKCUc3JO70wN1C1FR99Ws6x10JS/vmzoBeXnAX0YFcdverDiUvZnp
vHPBhfh0Qzx8+Pgu5+P9g2MUt0Vjpks40WeymWplLY5bYM8bSp8t0I65GbyLS4/1mwp0UvuKUpeT
0m+Q39BvSD1wQAGazy8g0ak/g7Q5a+e4z1d5qWFTjeNNMnDUfR+UbJoDSQQ/AL21Atyfzf0SfVj1
1/kxOdrrtLFfFvWPks/Pu2HHRBYjOMtmyE/V4Ai07vPSVvlbMRhAlJqp2SEqLCULehfwxF+Q6p3K
j/NYJDzl1TenlYCCYAM3JrOPTr9uNehc01fkFJ/r0JvNfV4cyDu1SNtsH9DqJJ6htH3jXfzFdRU2
B9KGeZn9AHOCgu9Pt8Zybcfkc0wt9/3SG7k05bT7k0s9rUOMJI+IGq24hyhz9ryugwwrb711cuAF
L+jKWaqjz7LT17YuA2IHNgK/W/nKFh/d8kMqB5fkUTcb3LQB0E4Cfqp06TOE5/uolKPkXdKtDkHM
5njfdiUCDAx3bIpb2iFDexWjG2URRuy22MHTTR24hR77FFI0AoAsOWfQnvsu7lalMyCjBIMFXfKO
Hxig2wHXxqLFK9viWXt/iliAbW9fTgpIDBI7R606Ij9+zspEYd01ZQrH9YirMPVPW7kH4iuPbH04
rEysw97pvyQceHHhELFl9eSasKNC0Bl1XBv5qhVmX8w9NHky1/kF2zy2H/JNVkwSLoJCOFUfYKg5
xTw3QN7GPtTKqkg+9fSDr1TQJdctfWYSLneEvr9Le+dmyred1vTKdzbTh3xqe8J8coQlo/DmYlQh
CFyWh77DbNcJII1JKNxtgbjdzOIICNzrHRO4U1rhEaiSxtQ0RbzgHNEp8YQpamcXhPGmtEURGzf6
71c/uIUXN3d1UGJ3RATWG9o4PAvKlZ2O6eXZGD6tMBRiMZOXoifoo2FomOZ4gbYHlsaSY+g0tTAH
wSPHyalpBRIC1cDiFF7JYZSmZRwAXYjw8sBVq5CMn12Bd/rXnvBiJ3a8Gu+X5k77fpJ0tqYS78Gy
cihFb/MblyiO1GYfSpXDKlJ0yQHNKxpxYns1dB4DuH52SnNbeeHejUyMMeTtNVrWzGgv5fel3yq+
QNqnSHb+8+mxztxCwHlJNLjSK3hUvJcN0MROQsLxdi0Fta9woA180kNHX5WvNKvpsk91XxLVSttW
5VLfRYmxUVGOWegftB87oRPbVROwO08z9o4+Pus5fT61OZWL+n0G1My5BNNOo1g54CnAH+MkDLtQ
EDjPmHtNaFoL43u0YHqHPD3MbS8j97Ao6DmwMTTVr28EGZPs1xu2RRhAVAJuXwb3Piwx/dWMjxIa
xc3QB1IqQbaNGiQUcbbrDek3eCXMhLancJgogHg7+MubTNYPoJFk1o0abkPliazTv4UoTyBZXTIj
5Jngo58f5u6ms+ZkM8dBiBvT2UF6C98dsn/qxgLdyn2oWkAGHRBkNvmtVfuLFmxZPOxzZrr2CmBj
Ntj04rRjEikLpodXjrPU6/6b1vZM6iakc4Zf5uZeeJtyH5AeHNAGgqnBrqpBrhC6ciSjf2aB+Th7
mF7WORVgJnEu7w4zR1rTKudNqt5da25SnBgK2Bht3iLMXkcSRDCHPg28ED6izeSCIcltFgz8HtnB
jXwGpoUEvFu7fT/ZVSJgk+QtfSyZ2fY1pClMClJn31Uq13xoaUW53J02wgkSTa8T31Hk0Wd7/2FP
w7G0A5pzOEobpw4qFFMZwFZh87744i5TAHrSZHW90QYF+TuRAc9THO5OPHUcNU6Xrkq3mpybrnTX
hqIgJoqzwaILrGL6p4ykXalR0kdFH9EQsb9li5u3Mv1zw0DGlK9Fc5gqYsAyxRlEc3lLIxFzyTQT
K4W5c/bn3yGmCnbLTcW4OhQOpDPz7/Vx1bwEJDVrgX2Cwd6AA1Ei8ngagBpqu+oNEJDeyZbiG5LW
mzkyfD0CBx61zuqSd8OJIjN4Uaf6C/NInbv9oCjukuhjtXEgF8KJ4660qfJkwhq6LezJp9qaklFh
THJvwFu/5wVZKJJTMbe8ToXjP3UmH7HHE3txCjjgX15BdTQmXrt2tEKy/sH5VK501bfi5amPXy3t
uf2f+Vtlavt0ZfBroB79zwODifnw7BM6T8CFZUb0B3YHG33M8jLNxIsAWJaPoTuP+aRJ+XppuNpB
t6d1KdL5DqYoQxcBtUKdrRcTa6pRo72wYkw9KJeWtaCJY4BinGzgzS2qjYlBxsTw6UxeOPTTWK30
PuU6S+DHVJ2/71cEWvDvcllWFNFCYVUP5UrBXPrBHYOh9AFHhpSgbg+Oq34ccaDm8JMfjABL4JyA
rR3MR5js9GjxcETMbKz4Vz7o6iuciS5HXtpw15loIK3eHGy3v4u5ouT5fgONoh9Yj+MU6WG+YEHy
bHIWP3tiPbdPaGbhGArrdpBly22e7y5iUEvaDX6J6a1hGVSYQc/7Pvh3RqAjZOEN+sRheonx9Ifa
2xxL9r9rBQpfnDlOc6qDr1fn9idRRbZgtZiEUw6uCQKXfDyCliiVZvjVYFhLUC21DL19GBlHJ6rg
dFFWI9FfLkzqaBuj/Cf1bHioeOz5jGRqOKIhncEqe+aEywBp8/vaJ+NEW7adBsFH17eBqViZKuEu
YV+UPyh9vZFY3wF8T//nZ5AAPtsU8q+XvnMGDpgKb25hxMFGFimKTmewxTCpIIO5lGVr0JL1JErW
E/coubXrHxguKN2ALoFrQ99jpfeL9aRGtjRdyyOzdG0AtTnVF+9uk9gXht1TFfPmuPhfL0tUV88J
wcpV866IC/HcTTfYWrb6I07b+jFrLhT3HZAEiYabqFFYUHWBmnjQnM3mpeUjMfoVJsnYkm98uzQl
U1eWqoyq3NB5JNceIiDUKw8GgpuDyUZ4QOE9aOQuYHmvdFW6Ra20h+KBJwmCxiBNcEnYonZK0GXP
r2/MnTHlrXC+HKYCK3Hgev1Ltzx+ZpieDyyIe035ZDxbq+YTY7Q50fSJo0n4i/CYXFKaHy8xlgVA
DHMPBJtTBubuazAxDwNLZBzmSeIvnhHLkMAQ7Fs+EgO4T4vDgsMrbODLQDCojsdjeQEytpygNFG4
0wtzilCoq2OpmJ7PUYC3XBnOONjh1P9D4iN4QWzHn2vaARr1lwkdB2TjIHT3oaPAnkukQUJno/2j
HSKC9Vw2qf/rwqqXkyVoziELqnG9jsbeEQZeHtINNPKZ6mBmnxtPFCj1uc+dFGS5miR1K9GjSYoh
4mQVvVPmJgXMxIeJoG5DrcZeFVOBTX24rAa9Ww29+2MHu4jhAXc/BcxZc6AoVG0ygyBsqLT9vMeJ
NS63Wz15RlWEzUVKkxoZliLAFWnMdv7Efyi6Vhfgm0BEswxCzt69Cnk4EmLqYkhaT2rXPJu8YOl8
BFGGyysngvl3fPLTbEAa2PQRpEb7f83lUMVhxC0F7S2wDvC87BovV9AiXZ2nZcP0LHGENp1vNPgx
AaFogwy/yi//rCbFIfV80Cd9ntWoLzRU6jkOS3zFdCg+lI4DrnQCWNhHISM5ZNVHhvzXddkeaMmc
ZEZrvZHQCmwZDm8wcrREOAlfe84mzmY2waTyIcFkLkGfl2B1t+lG9yS+47ZDXdZm9q78TGsgMm6W
ezTctvAkahDtCBC0APOG9NOf+rbe7q30WgC+R2haRg24pltcjVUDDyySut9feZtJoudDUixT6P6R
USQJ152sQWRhSPdqouPiZ0L4f0kBAkTm6LBbkGl9GG8YVQLQbv57Jh2s5c7pOP1vk321TQf5hsDw
xsf39fCjnORS0IgJV6bNppGHnhMIw76TKCK/rfsYtPe2fq1hhWdqw47N9HklsAgxs0Wf9K9bGivM
ijajWmP/sAGA0y2dcfTtMwCxaDK9CR4vZQCMyGyrql/N2j1GoCyIy5vYYH9CGwooz/LdTSJufaZb
8RorwiPtXekGGjkfORyno47zDZba48k7ho7mRwkC7raGuGBfSYkVsEy9EQOSm+hKNScwxrbZE6p9
Bqe5XQU6wSwPKw+dilvhj4y6jsMbm7+VEFhmA+6R1yqLU5NqFt85oaCGitmjA2+eChdaJ1t2XTcb
VtCL8eRkgjTEEnQ8XGz1W0qU6PyqzEvDgibDOOX/2HL39S7xzpAOuDnpHYvwhuj4Pulf11M46TVR
sKIFpXqh6ug6bMBDsozZcPYzAjErUC2klDHNo9rSKqQ/YBxjGE1SJO9xAGSMxB3IB6lbVhDT83An
hAxQNHSgrK4KBiarfQPs3iAMKLzkX0CudXroLinDRdxES2uDK6VUwB8EagG7QTxj6eTeJdkwvYaZ
FFNo/AKTUmi+1bTe0QjkUgOuiGw4gjWcadqKM73lO0FbRRM0J6gjfXKtuDqahkje7nie75eE6KZg
aBdHy9PNR1/Mvxe36jz8qmDistuiT539vG2Qisub9UxIEd+b6qFYC330HpdcQokBrxl6ZC6hgEuk
2aTsevHYkoe3LkQQ/ty9Us0tqkxAIVz/mdb6saAvjtUgAxnTb2Qgz2WMeAG+fAVAFiYA+xzgzEB7
0ZmRiquwAtK8wNBYofcUqNW4GFK5kMfkGOqI/LJo6EXXsrHC6kXq4Kd0sWNSQeUX0hzlLXrq2J30
ZgaRguyM9CTjvd4qdEEPf1far4EdVjE+8RzMK10v/Um6AN+FWjwPbTGJm7Pqq0RT65NjPuatGaQV
AXUi6axMZfbGx8qIFAXh47/Cd/ZU8oN9V4Lja7GGjnNsM3Iv9+hc/PYUI0mG3e/MRVUu9qu0Xtkb
F6BQDCdqIDdQxw+jtOgj5IruIOFaUJ2nkaZKfLaNWLm0xDsrIGWYEYYD75iukxGUcXjA+1pOAbnm
fGe4BxLKumJTNJZ2Zy4/RgptuZylY3Vr63CCdGH3gvWGE5xO5TDW9YVDk1EOLu96Z9TQ3olIiZFM
tmrX4SgdIQ7bZrwgELoXuwjyGUVBIds7jXiBNB21LlfCKbh7eJOo4PY7HRdllfEKFwrdKxHNfUoC
m9f0iikU/x5OPXRDyYlXsDNkJsM0fK3OgIX8eqU+TVXwQ8/ATqD28Dt64MaRtgIt78W17kM1Rz0K
B2Q1wwvdLSMJodidPdIJx89mxmVJSQLroBO8RbCMYFNGW51U6BX0H+tkYqAtjSbh9fTKly/YcAvz
HyARlBY4tp6mt16sm3Z23VA9Ub6G3aUopI/U2GYwWuePb/lSFovWJDpPJrFE75Svq5C93keUb3gW
3XW913NwN3uyyQhYuSWSwYAbLgjS3hB0omiFk/SrhOgTpRM26RZZuoOnzEsbn2eEceUfhy5wce06
LegSQg4MqRGxSUNx50p+flMuoiqg85GLuQaehTovdo9j71mWMoAoB3f65IRI+r0t2W1VnEIsfIot
hYKxJB9sCvlK//h3g/pA+VtB6LuNfASE4QBjTf36fpbkisDmRvATmTAjfDQD+VYq/oapmv3rmdTz
nF0pQB5TWeFAF8cqVclFPWr5kTcQ3owtaXTArUm3YQcYqT54P7QuSHWcz9Ij8MyqzTP6HBRFqsZR
abXAaca+jEFyP9b4pxJRBJHm2T53Jpu5rrQIAJJWTJ0es3147mdfFgvzgVIfa89aoQI3xlQgFMLR
oMBG/Pj6MYnQUFFGSPLKxSa3eJeq5hrEYsmkQ/8Y+YgsKoMhfG9CFPIlPmKJNy5hog8pV8L405/v
5vkJ3N0efmnOVl4/21/oQvwUGgwXnuXTBLRuZzPkXig3yNlAnzFYp/3FQ6qpX/jPjAc/rzoPJjYs
PK2jmd87009gd3TlCrbCakcMyZi4hQVDOpCCk9INNZZ20SYhRj4YUiT23Zga2LTzCjFy1HjYedTS
bdUod8bJtTQ1vWKL9S0tZHrFiKDV3mTKAaX4n2Miuu1fSvkCX2Q4xxtsp7QCIinulKlU4+3QD41J
M2gYh07s5O791IsnTyWX8HLcKr+W00SDyHRZ78J1uqYoxAETJ7DzqqhyYgpqEbBsfI5KUdDJS1Zo
gbVDKfCCUA8v+8sFzDpuFIk/D4b6I7fPoIW6Ba9OWKL+5jW0sJI8oEFtHiAfYBhjNsX9Axr9d33e
ZcspDi0zt8YW2iekwKwG0avnTQ66i8a08htaQohU1GBYIUTFLTiZ6CrT2HqV1utvYPQGEZG0oyHj
JOCRJBPud1IhFMnlNzfvx5iUyI8W7IWBmXtXfvxs1Lz4bM6Vr/ZV8ooLUt5+Dim0cOGGEfel1iSh
966jKQwfnJMPe3Je0/H/MUsNVNNcwUuxPt4wKIk3THVEBFtmaFQf26BQp8xDhAE5PXEF7VhUwHVD
c4847AJL1KtMr4U+LB8qgDTCdiiFjttaCbDVKQzDLNWnjuj5PUGUiIPrPXNEajxjesZOOjMCB3jH
nYCRRD2mEu13OOPROIYuX2/8k7jLvfKF2tHNOw4cjVCxoETtjQbaKIQXK3A5GSlbyVat1LM2FQLk
gl/qP6eQlX5EioAxjOOukNVIjGfQ1qeQ+5EPvy0E4yi48AfcbIWwjiTyS5yl4MfCHbTcI/ePobyv
igCtubfmf9n8690yNZY9bVmQa3I6ELlDn7TsO+43mA02bUP6Xs555Hm5UZzBXk3yFKCB3bUaOF6b
ISpkohIyVqKl9plIpoplaQEg4hh3FxCxCsnwtdCd4C6psAH8/lyIOjTOiRv8wd/f79P+jAh8MQLs
5kEDR9Mphs4ioY5lHBFFZimjyAQVir3go8TWP2WHZV3OXunLrCd/Un0eV5WNdnRmwTFHVlEBeZqe
nkuJzWxjQ4q5Zpac7Ux/zyrPjCE8+AduHMv+oV8/WtbvlApM3bNYcGTVjbNNza+z26yW5IQnFkIq
lzaCpN0D0M9xaeHnc3yl8Q3V+t/yo4pJ7wbvlDQjyFIUe49w3ziyPJbVDlWRJodmYjMhEQVryOZa
fpNs3U3paUGUxEWfRxvupRE9o5WjqRcYaGfLlk1hOm/Vz543Isn2qG0+nGhJvHZ3ElV396OtUrP9
ZAizRozu7uDtltZJI+VhI5pEtXR6j5IAiTe3jiLfhJFPIM2UlaTcPqtNwiB710z5VVyQZNBv0KGA
2VBq238LV3D1+4VoIemPs3I0k0b7SOek3isSnjMtQQqe/B5ckxIiBCv6nOWwqw5g05dSSvwlhfrW
n17GIhv7/6B6byx3NdE27YnlIHPNK3fQUQeN4MEHxCjVluG2jI5EGKgd6nlEcpuCuJVMR3LKBz/y
zOMMj+5h8rLRyLeS5/lzVskg8BHxtTocvPuT9nPdLiHJC7HEW3o3bwX6LiYg81rBh809XygTseIG
tLA60eusztqkC+WXcq37Ethm/04+3cZvfGZUvMn9MW7/q8gBvrBMkrPzA7dK/g4hrcYn55B2FBug
YxO43lnQWsZ+mZxCMVCnm+fBhmiVwpYUb1S2B12LpRljikrVxpbuXPJiL8rxkulrMqD+RIi+J5jY
Rd3Kva4owv11BK4Y8xgG9c5UeZrU66DzgMwHaFaveeZ5vnTAHkN8WVvvKziuWzBpi4dUr7QzDwXK
yBjZZgOQ0XFcPHgdVspD9BNsZAY95RifiPuRjn0GwbsRepLfWNeE/pTJG375rxnp1vJgrOIct2iO
suOTsMra7NtScHsY3dJ5xbEBq5UgAEZnCBMzyZtXR60DxsGV9hX3PDCqLrN/SUq4+PbsZ7WdtF7S
4XGvV6yB32EjZGHjpYwukyz7Teu7IsxiGFtGF/wZRVU+WThSYyf3JmeXwvJQoalqDiwz96r6UovA
S5CbQDHKht2xnoWqHuH9PYl2wZOsoejMzwIpN4eibSeF8wkHXoGATGdoTfJCnH20KzbpjvZMAX3y
Vm1uf7w/HdLn3nOPRa2Htx806Ln2cpFn3CUfIfhlNP9ZrLxmRs7oJNQLpbHjqZFUtT8HR18Xr5hj
dOrvk0HjgoSS03PqT6AgSao4/eB0fbLn09SXaBOYzGAL0kzo2J2R+gxUr8sLOFBDRBG76KGLu8DM
IPBALt9jMQut7/9drz7M95xUZ3lTFYIVnJAbJsWHzamgtVU4bbOM+baU6bW4oXq4JReVoEiorCpo
fIAjGyackgi1PkWlJLsOmz8xyqQ71Ak/OiY+Y+Dbs/wL4POQqhbvXzkeD2vMS12s3YFCX5Swt/pb
CJoTz+o/SgDvCl9LFr0Z0FCyFjV6CPM8X3QKQyBZe0X/sAmZsP9VtHlFK8P9BJfvuDo5y1962+uT
ld6LNpXexhPiTKZKXdRX2EzZEt5hWO5bko6PBCN+cRh6OENuVZZLlwYZeLVEqOT0TuGuAFpoUQ1u
uja9KLH2sQYz0DBV2F2nN4YAnIiJIlnFbuoCjLwnq/TAxFPvsqbD+lVc5U+TBJZgyioQH0K6+Wiw
LHw6/0giKejpPJWi+FMmX0ewn5YRw1wOHWj4+lsJsBFV8i3pSZQixoW3igCz8vj0LPtzK+Sz7R8/
uVZISFJXO2ZwU2Jzz3uzmoftKBmvXLAAVTb5KSV73qevaUfWmXrkCwqJ478CQAIyBX5fjjXIpWNR
3FWA5FKYYUXR/PvcskBzYM56drcmhPHU+wgjC3nVc1u7G18Azd95I2gWL/vRLAanCFN2mn8F6h17
IDDuN1GAH0W34JZQBVDHLZ7zaU5JVtmyVns2Eqbv0itLvVH9y1QYyrbzpMHvAp3R4WIQb1nLe92Z
nXdec6rUzErCpxLLSe7hjWfiyy+NGuXbxYek0BbIbTtM7N69ltvgXrhdC56Wzy7z0LG+SHPoop5u
gAkApPR05B19dPkueGE+ruu8kkGgiobCPfmBGWrw7OBPZ9JmXDTcMRhPZmIqFTKLlRkjQYyxbT03
hhu8J2uKMd1aTpb57a/SBSm1R9DiHfUzNxElK0EwQgXJDjav2ojDH7lMBXyJRfM8wdsHn64FeTAK
OiBLdsTpcWK7fG4S5da/Iwgy+gTRlW2UgaazQz/CjluyU9Bixkdf0ei8KoJPzmF85+sHZhvMlllP
IMNd7H7RQ8gzn36JnFKQHdsSLs8W/bql3+deF8cRzfEjeC6LcHQr/O93mp51rVT1jCmqd8YZA61u
f3YZPR/D4830s08DtDvIvWFD03K/elFoIv7Q/s2kAxCT+dOjKsOhWOYGnqxI+MagIzCzW55D45lQ
hr6H5FUSC9NR2AJv6HLyVaDxNkzJg6PKOFwGB41nbMKynuv+JouytcnQwx5FpozRrLrnLGgaGn/J
lSEaaOQMep6UUUvFw82q0fGtSndIJXl9UMHoQInbfcXpXKU+hyruMd2PkgDMLk+ihPx86iINwqIl
9E1OsRdSEdn06FjZEO8sQBOPvP1X5X+/CnfQ6/UwseIrV2SrQVSWUAWBWAOiWwMqhcnmr5Y4xs38
3Hp5gTwTrk73EOOhMbQNnYiYe9L6rLE89bTgJ351mTTdl2O2xpdMEOfVOa3nZiENgE7imeo5Qaev
CFJxtv31gHNkdCgGo3i6Z5Vm4M2qCPBUcJ5bMGQfzHwCRZgg1RkSPhp/S+VFGaDFwF3w/wla0vl1
yDEBO9FIG/ObfiVaPvNjmGC4jQjJCixng108Y7hTQ4CWkqBenrP/Q5UyfYARx6B/+p2n7O9WwZED
MyBJbi0HU3yNKcrR30EbZiQFBJfBfIkNUFBw7qIUCYg644xfS9pl37ukF211eMjk9W00o0TPKwrl
M9bjF6vbbV064IGqkZcTvCL+6IEspHlGMJ1iOe5xAPuJ5F4Q2Hlqn83aPIPaYkHasU7K8nOQJjwh
TcLdYZvcvmM1Hq2fV3OvId3AeBgTDUM9zC73qZyCCQGBRSWuq7KtTvnZXqcxCBHxCAyfEKqA+MXc
zOM4t1paYcQiSyqKUPgOAoeIH0rsmWlmTmXcZ1gkOF8UvpJM7R7ZQFhG3DXNKUQipH3qXqvbv+ik
/OaDicsE/E5/aLdzh6yPbjDs01zgAo5ocDlmrRa5llbYcCGaUNqT7ne1cWHVcustw+KONiZyz/ts
IBE5R9BdXkZDsGk8L+FJvLA0m1DNr9Tq2qvak+/1MMDTHoOjosIAXFe8IvXs3AyrleqG8P7ST4ZC
XfmxpVevPOWOc+SLXOOPq2RHHOMOfW4NhB52qOI5WmpUjvjIiS3Xxjl1rXhSlSckgWOtZOE60+Ba
XnbfHLx+hR5hmySzF3HHv5PGBX9WWVUcuPvQNXcRcJUrpJ0DxK7wr/hVAeWxEIqGki16iIHpvU5k
M5CIl++MzXxyi31RPcT/3mk7JJ8nE/mgPlTXipIbWyDA16tWfPoRNeI/49TM9C65k5ZhfLsxc5T+
EeUoc9+2viERI9zNLX1qRKDlXQT+krMeJ5Zu6uMScDjjG/c83vZ7krWjuwBaWrh9D4qTH42Fzsa2
RrHKFHyjTUkc++XNZHO17wHu3f9WIJVlSijNjzxu+3o2GhJigGRjb/cxKzue3Hvyfcrl4JM2HZsp
Bpn1iKord0k2/ED5JEjz3MjsazlQQOAzheZVJYfgpumwLVyFY5x6zHG8lpOdpVwSLfi9i2JmQDar
iw1MzpQ4fBQbkGn+FtCsZhg2eJtoiSsuzml9s4vKXI1Q8VjF0wCBDLqMT/GFjexjgZZ8MO8cS1ZV
cd+4/+w180e0u9WXtYqhuZmpvchIRElzHiy4JU7QUGSTErloFLMQK37M7d2aGTp4px+bFQ97m6Af
/D781GlIH7PXojaz0u8PukylmbyR4EwH8ov08LytRoUkea5k1ENBo+xq3gmXv4C7kISbh8vXCgL2
AVjdoeq5mIvsa9zCum41dndAsRlfABjC6yWZZQt292Yckm/DLMavMHTj68VjB+UXeelflf6GeG0i
or6F46+bnSc6PeOtMsnHsxaSk9cYZKY8O051Iv2xQVg7Us76TA8TLFXRDCCdPVWDcosCQQ0I/wH1
j7+FL2yMUNGQCaAVHXkh1ALc7/DR9xLIXsyII7lPovH8INmbqywFxlh9p4QtXLBezDyzB/BNYima
npn0au6p0TIRYQTh/h4d3/CTzE6/lIgN0nMF4zB+3H+KJjjDvl9yQyaRqe/8LK3K9ozSd1cdtCZm
zmlwjmYpz9ua+kTmtvPokfLvHGZP06FmtJAxA4m2rwSmHC4dSzL/9BQGst92i9+n9o6oHFdmnYi+
u8IjAmRkucORq3dTrRsSfEz+NkaYCr20TZSwy5bPpKdrWhSQwue0mLmy3EpP1JTLt6S9dpHvt8po
dlfptEoqWpnwZ1lJI0dTtg+eZcPTRilNAvPzaEYcKVtFDPkFotWdPyz4oINaNC6/wbFi2pUwoBBE
nUVPGE+k6ggXZek9jeZe+PXfgoufz8BJr3/cWBy9UzE9caFTWah5t9esi8/ze1P7lsYIx1om9HF0
RKItvyoV1VKNRQAgyDISshAXvsU85LUV67Z3aSnS6tn08IQDd9RbgQiRf6lV1WMUTJdrhEC404gJ
stFXaBw95j/2JZ5F77/qoLpicnm+KCtKvhmkfrOQPGcwIN6MdG/cCrIN3HLvl6wMeOoaK7doa54c
y3BXw/nu4lEof0Rzl3c+SNPNDWD4FRydpuByrY2/v+pr7aSx+E490bXLJi7vzSgeie/Ic2AqftMk
gDO8kp7iE5tDZ9SAkCaBlJbEWS2ohos3ON0wsLJw7G7mCjwxa4gODj2ptBwvI/pMAjfasZcwthmV
561CCfh4WWgTAwHtvv/kik14vNWYEvHqE0kTxjg5L25mG3mUECfFGXQnLpTW4ny3BQQ3i0o1O4Nk
yaG3V1/s+u1WtNh27TV2zbqXDr9sP3WyXWYQnEmnIuDwWLhBDwPkeRHS2qpZNMvcsEUlpxVQutny
lmel11RwRld1JH5Gqtbt8b5ozP/IemtPfcUzJv0Zxlo4zUszT+xdR+XLbdYwDZy1hOqnZ+2j6zxh
7/OcwknQCOxbSpRII5cZl+KpihjTBFUuv5AmKy5lsj/VvrkqHBMGnwOA3QO7TC8ZBfTogYhFCq7U
p1h1Rz+iaJ2aeLWjemERz8jssvL8ATe5aUxRubhdbwiCkaZFKTGfLrha6mHaLm9J0At/kiesh9Zo
Nbd2QtRNknanxXf6cJWijOZfNNbIzp9Pkgm7T6wcF1Y0NC00G2IuiEygA7RCtxYZxmwcpsDsIQJG
MhVv8hpjrUmOxdQh9Kv+UMvL5E5+Bv4vrsfazqZP6m0sJAJ9rntWZ/eRg+da8jXP+DePaUwDWyVG
pNl53aVWSCbT5aSf3JCYZFCkY+MSI1WWiTMOsQee88/cqO8ny9M/ThQ3CxPmvfjkHmHmwg0j3JmF
qFhpTv6NGEeWky+zEej45Q0PEQbR8eBD/zO1Awz8Rmzo0Jk+nUjoOs9G78jVCfn12uwy35nuHIHd
TBRr6co9My0Ucp715qKXr5PWSEm6UFqT0eUQx+UnH8kDIDSGhW58O4hAn/9AuVf8WQ2+ZeyjiQxj
jxyLjxBCe+vBr3TBONtgaD7aJAXW1YA30y9ON7qxbXvX7W4uU1EcEmIQhSp4CJx1NvUY8lyddOcP
wsBFrpJ2/A5+lXYLyiyTrw23lFGih45xh+7OKGL4FNDsxgWgaFi1/vhPCwe6FVL55VldXxPrxTdk
x2+zYpR4QKyXxSMqQiI6ZAxHzgN1vQJKPBHLcASzJgaPUY3WlKy++LRq67JI49XjrsJAYoup+vCo
lsdW9Jt4WDmzUqrGgs3tGokPbvf5CEhVg5eyJR7MwuraoxL0h4tk5PTdvPyCMn0yiddhiX3UcrYy
pnwOrsNtm+TwUy5Qz85jk9ORAt68g2EDS1pClRD7FraCGyXomr6LPf8yzOQ/Cfq6AyasLTr73EQd
9DPeOekJbo/6qqbkTb8s6dlpq3hXJTtWXv8O8yMTEQ1yw934JKhwoDyoWBGJ7mJj9B/YW+zzLbOL
0WRmjXn7MRvTU4fXaIr3YnPwHpVRIDccThN46mmQqyDIEg0RiDNhtRQTUti1lS0Xs/DRXnbt8LJW
lj8Cx4o/Jja4N5W9uLpkWAYN0Zss//DiEZJmGjhfMJ1J17kVLUawhu0ID9Bf00ginqP8aO463Yl6
aIaBaqk4Cv9EFv43euV3ObvAjYOsLaZuFzrNo4k+Th6t1gtiQVWH+4MpRT2PqefwQ96OV2vVLWtk
8NNz8HCwgBcLSwA9NX4tLiDQrGd8UF1x39KuCe0/7yeAOEFWpQuzvZACyMNfd28/u+YcrUYd54kd
8zv3va8Wyzj0HhAiWosIvKuZCmsF95WSL5NpErwt3ogeJ0syc7gVgh0bKDBBDG5y2U+Q9UC64jtJ
cYWR/j2an6BZkI6sFbKAgzYWDNEdaAsQADIF/LmbaBvPzZr5A6fs6OrpVeGmaLET8/wNMs2MKNI3
1M7FRKCsmBxKqbi1JcOtYk67JMf9aDOt5hufL7iwXj+hW7mbs/7IeZuWNp7zhh77Q4451BoEyG/M
iP+aNLxJGNQx+owhwjeB1AciZ4dhICETOhvfMrziuNjnCvx+L1foKgrRy8domQ5m2Wg8PzribhXe
TLpvDX/9sWBiNbK+Uv9kKf8A0TLK9n7rbdnBl81L4QQqDi0xg3KwzUQwx2EVxxcNTEucc4xhEX2f
JcKlfWtbsCA/XKNTdu+mWtSO3gTv4ei/2Zz+hLuZW9EtsHLggK4CvGGVYRnNCNbuwQ+oMZ8K25q6
9Px42eAl5PTw43ug/qFzt1OuKnEyGtfCyGVjQfYqcCAyxgdjuoNEYDikAcIewyNkZcmYbIm9NNO/
1LdGTWx6phcfT9IIs1dRyNBFsxhTIH1p7GEDS+ioJIh97eKUCtUjzqnu0/7nIF/kJRw78gNk23Mj
bjUXUjhrifAnvWz4SEYseWLJi6sdUkFfSLayr3FfsgoedBeAqQXgf4xSqFst1raVlKmi23W6TJVB
6e73VABHsQwGAO1JiP92q7IiIdV/F6vp0Op4u5UrWTQ3R7KqzVnv6QnkYKQYiHNOB77n7HdCKFcv
pxNwX+xedUMS0g0l0hCYyvXpvIJLcy1e9UCkb6/bIK1KVAQShPBfACHDdsTCvFuD9RO84UyeXgZs
PwH6LXM6nTWS62xB8PyIDH/f7GC21OUqh/d5zyduwv5IRyGoV/+9IMv9LT2ZxXpN4Ks9tLXWyjSU
2yvbWUd9DpwjmDso6/cHfUgEwX6HuhC2Z6HLAzsxaZV46uqQleVEzaHOPj+zzEIvEko7Zj3EYUDP
4hsdO28MoXjI8XoaG5QBI5ux23cEMhjIRUADQSTdW7C4d4/MQvL7Ea5gXOuKvT66EGqEKQ03h9ne
6fztzdqC++ea5fsP9cL1oZCYlEDXNxUuxZjW1umMuJhh7BgZj32Ei2lp6TcUwPGfzFR1W5ZgwER8
2ThzSXcbFC+/j/dMHgGieLD6/s8IkskeME3lzSLtinoRUpW5iuNfnSqrEh/DVfTYkhsO6gsV42xr
d7t+NNIgBednT/QW6rjVAzIKmcvGKn2U/97Qa9V3FzFhdAKxk5dBEurYT7MFKZaEoQMtAZo82TsE
9y7Bsl4TZfrtSi7Lw+WFaikBrGIiKr6wTR/Ge/S3eNbTJz1969z+1Md1HXtOm+pxsskHotVI/FsG
hDmfqiZtLoVIK03GJbbaL3iUwf8tuuHgiy/oHIR74m93aNIjIAOab4evXgaPMGRnAbcEinIOTNt3
vSBprN05QxuMA8khxLO2LrY19+edHnvBRX5zooqetstuU8MiXs/7L63dEt9wp6BRvYg4v36lOdp1
U9qAlhJU5/VlU5iblZXPYCdidAtIf81nqSQEE75AHI9Nl1awrBY3+WXONKT7OwRqOUN7vHfcuexM
3bNMISDLTi/s9Cu8LfbVuGvMtoA/Qj/xTmLhE4DREix/ThEGqZxgh9zXUY5ZqzRC9pWu5Vn2HFSf
kx/DO9RPYHvi84g51zp3tg0I+tN2E7RDSRT2va5flOumzk89+IRx5k/+fwq0w5hLrLts2GYEZmq6
UdZ7b8fPRQLr+yd1Z412copxgivcovgWzwXaoyRSho2u91qTKrKyfgR0N0JFBmSriWzoe3IWYGqi
txHdJ1eEFw0rewSqgGifI3HQmq3XukbK12kW6YA96YmCthhQoUTCBzbVMU4ci9r/9VQOTUarf041
hTt3zuG1+McEPHzJQIej306lfbuq8UCZpsSWazXjQuU6KzrhP9MeY27s+DX9rCJbIQrMCUIC4R3z
vGpRbJzvnd68/yA20YxLhSjw/hTkAx+X4UXNLQ8RSazPsymBdCrobO7Dqhxdiu1QPHRBlggRRvVO
Y0YRTNz4oBw2mXM5jCrJ09Z6Ba6XrSzo/1jb79+ldvAQrVZt0A2VPV6aHULEJjPjwSNs9g1D9iNX
nI2hSPr6phU3qtsyOh4qGhYC2jPiRDE2LB7TQ5q+l6oPkchPC+LYqlqlNoCZAk81eB/ORjgru0jg
4NOC4eaaBbTKQMPOXD5OBaYBwEu5kgp8CUd8fR3ziJmEd/rELxpsjuib2QS4wbhQBMHh3tATeQyx
DR/uPlxumSfqe7KP2t1tq2TNUMYlDZmeSyr9LKMoGGb+u2SYTXg7VgqvQUJhnjDJO8IIDv4bOQkl
4JUpsauN3cJCQKok7fo/2GTdmJEIMSJUoZGQZcdBfzLcM0exdkajWXRIQmkhFbAOiQDu77sM03lX
LS3SeTuQJs3rwspN9bQc+0HHC2sXYj3F8TpWBqtbUqplBM7c5p+ONDsZpgd74NNcBYuzOhbLA6Jp
rw8u5oS+TqCaNWah7JfpXmNdhX5lAbNmdTStRyLlVzdAu6/d8zNluki75Y4Rv5VL2D8GGOws9oIX
ddTNoFy8cwrTOEcdrJBkguLjMlgEvBIAXlKI+CkzLew43Spcww10q/dHKBLHSHqMHTk4UViLHt1W
ANQvnigz6BT0RMs8VMI57JLUByEjKitDvcZBhtMsGd/Rvm/4wdVEH/gurGNgVRu3dGs7X4OBSlAw
J95NATEGqYNzwZmGerXuXFqauIfbaSQ2meICE3qvjAEDyQNqc/X2PUppejsQpO4+Xost7QkOoUeK
akHNkCLM1EqjnI9Fl7VSzPJ0exuMON/vy+LFvpRmm1UJL9/Xqba2yY7azO2oMlv/RTIVR9XSLesb
YKM+GR1/5p7AF+AkzFIASjBEiSScX9K095+PawC9n4H/DCGVGw764Vhshk+Q9zrB7zxIGionL+on
pqlwib8uaupCU63JTn2kc+U9vThbwaVpriYWe322QwDfdwsXJUwygz6JqVxV6CxMA41XnhYT0czi
xEmVCq/rzrfj+ifrC9IoViX124Cu65pTZsrVRgju4m7wzNWf+qnCfmrIx1P5p7FhGvbEhdAXc63I
oAJBOQGe4Au+94xo6fmvqwCA+f2lWgkJ+GAXK8etnEuJUZ68GiLI/k7WqhXSa83q4Ftceew6li40
0ar+0Zg3x6syZWY5V5FuCBcRgsrL+zjx9KMD/iqmcf7MBU3ibWMyfy6WkzVVek4TLwODmw+xZyKV
IgX1TN49HfZnhZ1La1U6QZX8u9H57K0/Bhh40KR1fWMgKFUtyT0QkfsgjcP6qv83qiMevDgEVmFp
Ke4b9dQ8HCQPC3Tb8azSNGaC0D3afAXQJnmVb44L1vYaBIdTLGyuppAEwN6gR7mTlwH5i2asGLKa
eYN6UF1VhcqTb0zsEvePwjOpkqsg9gPsf7kOXL8XgfP/eb7GxbH7cxtXpdk1MkxG9lOi2942vaij
JBFfGLGSZOn2mrJbl+ABPzFGpMTEvYiMAx9C2TCho+PiU1rr9gcJHvRXiFdGuvQQ5RMqN4/qLkfn
h8/E01RHcW9zA4AT9qbkM4fIQMSCR0B8ESFz5oknhJZyxGH8O2MDj8uSBQdt5614knrFd+axcYxV
vOUIjaLpyVnLYb9IBGVK7vqIyNzCermPGKkqzGmJGTyiqmhM5Od2iswZXyLwKcF22B9m/PBQ4y6H
vwE0j2tRjQseljd8iT3YsF2PRlgi96qeinr+uLTNDyVns2MJzhK61g0NdTjIq+IS8wO8nL5EQs7u
dvwoxfGGiPcODlHwhGYo74SX1LPvCxcBcf9gCQZZMyZmsTCNMwnT448uOxxXk7d1mAMsbc/M51Fs
bHCQP0Eo9i+xHza0sbnWhGUy6WiofmGwx5ZcCfmOrKAMTaJfpPeZ1GgO1/4ByaLyHRI0JRrUgUtK
gFd5QVEUj5q/v9ZYdu6jOtdnvRbKiS3VBlU5oMfJuAoP8zXavthauJJYHZb/JqzG8P2rQC5vOFDm
q19P+QW20EEWlAWK2b2hPX7j54HWIRfCNnQPEVUD+u6Hm/KII7Ir3gV9FBf1Am2HNAYnPqYCnzVb
q96kUXjOgUHn7ay1qwoSJcLTpHto56tfcoQnXwY5HjSZkTodj8TScKHJHAvLlbYpwylO6iOT49H4
FqkvbXwg+k5crJwAvFzC9oH7L6xTCOIjLEZd9dtEywg8JyG9d1nZadInOzk5tVJq0uRshXaDhjjW
900o1baJHY+ourZ86VIX+iaB8RbQAvjarcVv9usKaxGFrzPWwKGJgIoElBSskDwHXNcy1XE9wyjY
Era239omPoLN0GhaD8aFcepryjaZjxGwUr31F992H5a+AN/iffSoPIOxg697LHAC1s07o5x2dMJa
kNfvR5f2Pl9/KSgyf3dhEuuCNdD5+tHrVNfzwrf8Ui6Qcq5cTiFyhCy7lhIxlh6s0QPzVhT2ClrK
VB0LqGejh4QTkL88rjl2lHcXAHCPmQLao7TvvR7VwGb537DLylEqrRwNm8fe9IdQND1XGREaINaR
ZfFjOjpPjpMj9kuFlT/xnUcToZx0V/F/jeS3Gh1NpjOoG6JBdc0c6j6/TZhQUY+tcLnVPKrpu3O1
iG9At59DpT+ggaVGx6nSVYDQbWHlTx6xYHNVmcuRWPMc8jD+mwLaVK+51EidGPyeYgBi7kw68Etw
j+Pbi2wlQa5ju8wpatbHG2Ii61YcejhOdWLgFFU321ZvoP0m/Pc9sUaISRnSOc+PDaOkVbHGyLSK
i2JPuOZtGCvtpJA7YbfdX70VvS0naR2D89b6ZUK+SvxGf8iL3vH9opn9S63jHmF57Xw78mzFEoUA
MC4ewfX1dGXAOxhWNZ9t2PEr3utGXStEjmZZDSmTeuVFoB+aaKjI8Abn0AJ6p5UXe0WhEpkeRJCg
1HXjIjXY7/bySrKLC6Xn+Jin6/640YSKXlyTabOJwt6gCTOBlaxwVJcXatnky40iC3c9xdk87RdA
0/FO8EPYxhU5D3hVOSMyYL/N/EUY9TTQO0R/qWBsHE/9OlyKc31/FHaE8DDaWqP9jEwy+4ePhr1l
8coIyPo7wMRANO2PASVdKxOA4xRefZvBCDlHhh2YyXKXdWmP2oL7qj3pzBmwaQagQPBRNXaR/TB7
HWFU4Pk9jzj0XGu6OXdZvSQs2A3fNcGgVFUOrrVT+CxzTVys00cBo6CAfOZK2M282jzFaEDqUWX4
ilD+cpYanfhhlpkYX6T5TwAdb6ZqBRzEJ2r9WpuZZdwJF5lWLKyLU0bg+Si4OkXLMrs2hEqy5lPh
IPkMYwRQaV/hUoPqTAtwF++WVKqr2OwG5dtuF56nArSExATkRXS0zXCHmZYXry5EO2/IoMD9cK0d
4zTrOfI12UWEqgvYLAyEGXJmI/np35Dd5sTVF6EwAy6JNMK3j79c3GG+7S5oI8/mqf7qDTo6eCG8
ZCFV4brkNVCyA6FnBqZ1CM4MxSgOS8Y2eDSUeqhG9VKFIYB2hDN6Su6hIW55Z1ChTDtGDtHOkxcc
+HseRxxPbWPB6qf29of9nLD4gxNH1DvjRVfjmTgW8nwvJcNUo/9OxWAwjvbDuALR/cuhCVvIJfn5
7CyhZBV+mUgKYXLUQTT5P2Lo9DMfTFGmEh4e1Obpr7cOzE8Um0Eds0C2sHftHMb0SY0dhJqswWcy
UX6i+KWI6z13akLb7Q8VH6Y/sCnsFxCsNdhNwEpowMHJJUdES08MRq2MlPlwebStEysfpx8QvRfl
6N7scEwCXX+Fb7rDGHdrZJ+XCiExlUqT0+4C4GIjCp9L+fTDPRGhTssBGeWNRsN85V2PUyBW1Pvs
5wmbrJxaT4bJHrISRjFFGf4tEpz4uD17yUAbeUEnADxS0eH1yBXJhklzgziE2dEnQYOWq7+4Xeo2
Vg19duQW7yHCbPj6xlkmx+Cttj3B4VAYIAibivEI1vRtPOnlR/7uoKVgofwIFUaQankp/wND7HRd
e3yfTub7cppO5XJDrBhkgv0YhQ8e4aRC6UfoWpiinUeLTm2hx5fiXqIkSX/M5Q3hCljJjarSFGw/
T5K9uFjX9VSzKDIf//qct0li3l7UiNMko8aHOpQXu95WuJkeKRLirtaCDYFG5v7GhZjPpxtQivVz
V9b6WjZVNPK9uTrj7cx2LeDYYogCr/6LiIuYCUqSZuGFO/7W+t0WuhlkH4WnZCMr5Zi34jEVgN5U
XYqmf/4AgTLjYfsBpS3/yaaaEYsMt1UOAjlSi6IQtwK5c7cZWun/ELK99/NfbYg7RH/OYvnTN56b
Etpusdy8ho9zA/Pk9hOf17B4qWqbFVR4rIcTKc4m5EgQGPK30ScbKlaWeUpx2jVqF0hlJgPRv1YJ
adQgAVG/q55wQOdmwKfMlXq6+DmA4+ljTPnJipodcEfF5igfJpkHDUMUmvoxI+5CvaXH+DlVLyQv
VDvksB8iiz0JL1oDgGiq5/94g6c9JNgLIdsfsKZf3A3HZJuy6oSIKLuFM9C6IfuaowuYnJzspNfI
2oEseIhfdub9PHJOxEubb0FRZ3ltMEw5AjPDHstEfUVVzZMtDlus/y73xJc4gJkwMtoKUB6EJZM+
pkMoo/dZDMP0owoc9F2Nu0Yn2vW7VppcgOFqWiiPDMtKIr6s0/EbNgtv1hBraxXkILviQySj6edr
d78xWgbFdTjCSrLkv+lVMOKOxzt1HHUdZPK/QEUQr86svNR3VpakRbe+8sAmgI5ef5xR5XegA4kG
f233CyRlKVyc7XdJC4iq9xP0mMFhuWSYrRcv4rNIqsxF1LAvbZEhtecEzAJeqxWKy5Wy3d1wqR0A
Z5X7cPaanZR++B/LYGiUWHs9EapnyUSu7XCSL7FcAJWID71n5fIZ6gz65puj6ghpJYmGuwpr9Dgf
D5g0rAKf0apUD7kM8lY0iH8lREAZ5tkI1Ml22pZZRsSKYGOg1eIjdg/nq2km0o07YrpEfV+bGVAh
IPg10yQ0kTMKSrucu37ut2untvinND5heZmTqCSgwJQy/nR7gsV3fvKfRuKBgn5ZulWzLZ026EAs
tyc5jTJq8ydrN2wZE/hP+QB4hLhgIOsCfIc3jBN3AZMlNzy8nlk6muVAlNTvldXMBwcTLC3ZPJXp
BW93i7tXiTpv7Qw6k4HiaRxMLfFCv8WRLcqEwPcBI3FMcGTZEqwrnWV9IGI19OzRnHXX8e9+7rAM
93u+9332uF3lo9xm8+uu2zEuUU/VF8QPBiDqEw4x4p4chIrAKTXaHb1w5r1SvH99F8EZ0EF3Bjod
Ry1FIVLiXM791ulUePyjRgAOqHUa8qkzy7YDGEnFAPdv6rs6raGFLJ6WfkSagEraG/ywh/jBaHbK
/2ewBCp7zQmvDEvqyxPtL6iSUaodq9fsr2dS4mntVLpuSG4Za3jz2wWiwCVGIAy6SWKVCqb2nCTG
WpoNoX+TKp8tckxxMqAL1Rv/JmLG+AD0BUamUGIjJncGcWondshzGuLw1dHRnkgZwL5M0s32Eoj3
KOq+MCcVn2XvW05jpBjGJhbFn8IWUWz3EnlVLFuHO6HCdC/zYBhr9o/W/TibzF/CsZ1KS7TA4YW+
Vb2KYupDeVF7lqhbXZpcK/ED/O9nF6I4trsETLMOkrh5oF8ZSoG8z2t4cmgZZU66WbJ+ZPpr3LV7
mioat5R3/BGaiY7LxssDV9YXIYMf3VfoyXOSec6ItOdzeaxd6vpiEBlS6MGN8s/NaMDIfaOnZgd5
xXzK+WKw3/MK9k3zOJSUy6wlsS92Du0/EnNVBh82wZk/ATqC60YxAuj5NKdonaIhrjgmDiaAFIrA
ajw5K3sC8ixd02WBsB2oZi+VyOrybUn6MBx6BocyysuBm9dCSv4JJpBRmjC/j4rtViO1wvCGaVjn
ZKqCxdSMshZ03MhQhmSgeGupbJZpxmaQqKK7c2c+2Rxxkg333LkON5+F9VwqRQxO5rp+rY4cOs9H
aCxfq58fdmUL+/NZrTPVi17QFirgMxnWeaBUcSdI293CYP1At4qj+6PKvGE5qCBd+RJKR3QC5jVk
ssxfqTfWJiOMofUV2RMP2D0T66Cvp4e7P+aJmZZeVWC8o7X1L49VC/LB9w0f1LxhJCLrF5j7wPBz
4/J06dzdopRUb7UdF6d2cmQoJkbs6cPudvClhrsODE/tj6LzCun7HAAD5luA7iWrFL9h/dNKa9gQ
mDAYeaC7m6PuNqPVtchNtj+Tuhm52MSEHKkxa0Ref54/DXh1qT7GEGbOdi4pVJhbNjfBU/p6/yGI
ggoy2RQdBWDPrrVWFDDMYcdhlMV20LaN0tKxAt6cieUcy1aWbjSz4Hligb0UtkI3eXLhPdAQN3Ap
V3YbIRdmv2qUojAkFZGxVcXmJ71a/whou5N8MHGZB0tY/q0+d32V2p3ii6RZxVktuPQY8o8QOHh9
1WLvx77nUpGfk+5BNHxGsmjJn0fKOhp9nc1/FPpof+jUiUp5nB1wRB5SegdOZPvQXwq7U4WoRFHU
EbMMprMUuP2SJv3JoDr++8Eh6mqdmId3F9YDRM+IhEcnAzsIoBPcQ4HQ/lnvEQWOBwguTpAd8l2f
jk6PoIWNePu8EUzxxMB622HTmXFLYYAB2mgJU6UNjZZ0Sq+3n2ZNBiBLA6h4GbHXd/NoCZQjqWes
jsFTt2/ehmk0lQPUvHBSIc+jkcs6QcovP3vS2ocW1lmzZMY5mq2WvavruOMoh6/yPtXudK+CzxRo
bkzaUhp8J8KfdQPa4xTCqjKNXGPynlUSrdysfHO2tuKPdfoRxL+4UfZUBTz0N+cmAIpNf45V93mX
3szaHmo4u9CrlShn2UZzrvvRVnuhD2kxxoCHnjMCjDpixc4tGtGpM6Aa/rLpM2BJ3udTZYH9BFtp
bi/+gFDwUzE5ZhujywT5Id22dSK+s49cYuNOGW1VZ+xyeL2aPxyp/DeBg0iVM1eSfoF2YhOTv+jU
Pn94Bvg5naIRsEkiTZ0xGKTR12FqgY4GTuHMW0QhRCdwh5iRXh6Mj8WKPS9pQgq7SQCtauW076mh
zenhQh7eP8L/lHiUf8HDs6r8SrRteCv2wQfOKXGUmei9h8AWFm3Eppt2hqTlr9NvIGRhqjdfl8CS
P8PB5FUPmeGcDsGO5FJCBcYdK+RRqpwadYTt7gQUhMqchQf9OQ0m7H1Tjv4dJ4geq1C2IOa01F4E
zAe+woLsIbrZx6E3sXBLfJJJ/DhojiNlmsPUylg24Ue4Hzynu8cbJCJ+qpOWQWI9bjris3x9dspI
EoT19mraEF9XYy6qYQXKL+hYvtc4nWwsK5/CVXGFi7JZCEgjC4N0rNNnsMsXhU8ThCXJ43ahxc/i
WGBCRvRrtPdwqyGLLCl8pNRlaDqfjUnjyJlSD9mpU9jNraZxH0InN7VzblRgHECJhOBtTcwKdaS5
jFyKBGEAi5Us+YmSPGiAIDRDoy26Y8EITExzXhdHH37yvvZI/L0VcIbg+u6VHKLzcYnolQCIuBhe
o0ZhRRjr2Mui25o32Kqjk3thoRgZtTBTSxv1Olr2betqljKuNdlbwQXtRr50VhLtukp2sJO70lZL
kesM1et6pHwAbXF/donleI6ViHzz4IENb3LdKeiqGNak2riosEo5O8HDkqGm0im/pkWdX6SDrMIh
ITtR39KHB6mglOnGWH9K3XUeuCXwzOeVxWg+bhXNDfbq8ZiSNnMvRx4PNRLI4VL7aJ3/8YsnNowN
dgLKRX82q/pwJTq7NDmFgi0UGWPJvVdHrBSWptNkrsvCp3tcT+qtRc5wyfUYiTBLN2ErDKE4LydB
hFzj/QqAeWtYWwpvTw0oI5dIRNoe8luPl14baATUsC0JUwpRt/9ucsrsMN9FN+Xm24ZafkHf7qRY
T8Cn3TH5oprR6j5JyZzDogm0bhzjHBz5RpTXPsMyepiOOMnCEZKWYY0RhLem/7S4KFIAbSMKoBcY
ax9WrCcshPc7Sks+it2jOIF9efbREKVo2byIyiYFyJ0U5CWJbP/cZMaTfRqDrTCOH6bPCvcyp6WH
gav7dGBuhSRkrekYjFTDSg76YaRNcnybBEBsBLDisnNJCwtTkIdblT1y6ZW0r2ENdBRZyT0FIZD6
O4oGL9erUlTQKQPoEsFFvuFAmZyhiiUpl6+1pTCWnspOhHehEA0svygQvoUV7smHSBDNMmKsyU7u
L2Pf0cjvLrgF4bN2tfeo5eVs2TB1aoDjOZBFEh8MMs8i/V6hXZMjW7W1OxhqxdDuhUERAkXtBhjD
QYh6j8YTEyQvEISmjezG83a9/hBCJA+Fmx8tHh+Js/jBhvhjU3PDU+g5EueS0cYEJ8yat6I3S5VX
NzukNduxDys9Hx3/zc17OWJAjNASUoRr9nPCUAV+VLErKY89QPyKE8XtZW0RLDKr+0w0UN8CZ0Dz
KHhdjZuwQ8sam39b7N+BWlLgcXdsG39ExNM3txPAE0/11rRx5hBhUycU9rELUufZZPcb9nwZ4d5+
EARnozpsB/jZ7F96fxhMxtlDsjkDFY9j1/guBp5aA7jSdzKpQuJV2gWn0Ru+rtAA412aCzd8D/nn
9p3hILL0iGcxW/1S9ARcNTZhOkvPLuVlFuDsZjG0mFJoKG/TCXmXsRA9NJL6GF7DCQK7F5qO8hjm
PmzyWU6MJeYRX9Gmex8nEb2TccwFdW+nB7Jjs0Pk85CrZSLOxWRF9y6ixzkSouogu6vW8cKNqnEk
WXuFy66OhXajg3qppt09QmLKSsNEE8k6mghwh0Jf1bYhn2UZwmQ8GgoIofKILNYPwS+b9s0d4ZCL
2YibirXI+goKyTViKFS7nF5lwTDJ1uOiNrJSslkK8QoOrOrJ1zBhxs1vIJle95YDhNNRcIDGZf/X
ACk7YlCVejFmtTDmP7iiLg6+saj9nUhhm97Kl47ZKT+26mxk3ETFf3p5O+ouWq2N/L+73M/TIskU
i0uknmvyTxevB+AJiasnhi2nZp+jeylVe6iYQLF6bz173FahaFN0jJBt6lXrVx4mTeLjZKvbCEh3
Rucrpax34EawvFatkdkzgjIyB7giauGaEDjZs+ZrSNDerJYnLJoTHbHroL3ez+kFGfiM7NAlPRPl
L1WGXcW5Y6MUwQIkQbDYHIe7SA3xwC2DoIfLCU9H0TuzDte5UrxNf+CCwzH7evDxP+Mk7nz76h2V
xJ5h4oFJORv2Oz2Ejgbz6BcVRkv9ZoQlv9y8Yd15vutGjcXYxU3D9kXlu533e4htLSmP8ft1ofQq
GHAhlYwuJn0gzVUQXkxXH+OJTdHznfxmm0eUhG9SpK7yiia/gnMeyZlYgGNFBwzK0RDAkyq+7QpD
KiQLFzD6h8QL8c5yOSVw0cyhe5JceONO4yDWI/eilrcHpTiU730groO4+U6cRBzkOo0G+ey7k/Oy
VOXoVCJjDdtyEJV7PmiEW8i1tdr1OMg8GxRzvde2G+sMrQOdfR6pr5A7V6iXrvfG+Of0fR5S2hsK
NiX9YpTakE/UnPjFx54ECs/2/lf563eG91MWixBYFNR/6JlsKNmxxD3BeAph2hG7TY3bfN50Z0Yp
EOzNnxvapJJSj1teCcC3bCDEL3941GWnlJygqlUbxah4VM04lqaQza+ycC1H5MG6JNH6LN8GDwqo
OjmSob1HPJaDbNvwhBYBoPE5DpIe4g5Oi8vPl3h66ZFZwfAY49M1V+REVVDQlnlBRMpsxfcZd+NQ
jFJutLnTWUeW9wbz2sY4MYPWRuWbbp3482K0zPnikMLL6l2FzAcv+9JfZ6Fbmc4gk0g4RPWYz+l1
YrdRRsbtu4XoeTB6+Yoo6F4cgMXEJmRaTNGxSZhESigmsDRMTREGAz3qD5SIw4NZHTBHjmSc+B5A
3moGux+/rRum5sF21YjkRadT4ATDGjE4q1DOhBMctbk+4c8GXWpGv5IAzTkP7pRFoXAv2g57xRe7
COjvIKrqaC6pGoU5wpzVDW0ZhLtlWtDqTHxBWeauKr9SHYneKnfMnNSaEkF1R3aTi2LMx/6W2wfk
zKdLCyjFKIEgWY1k6JwgZjFjfTV1gIMDSofV9uoe4wkz4rsnkVQ9datP6ga975nnLTYYCW4/r5oR
nhdTPawJeKf+4iABkrWkRZ4XDGC570lDnw8S2dnsPZNqnD45DyYwMNe58NR6vgxcYCAZt+lODiSf
mWF7VYamAE9VwQbdV+blN1xStTuKp6KpsZHiOOvsdjLdZK1UyRWAjWEnS0IhThWXAgkBGJXKztJL
Q83FMh9jp3Cl9D7/k63f9EOMfd5u/nLOSS6qo4X9cqv3F9e/eDI3IvFDRrmg5+qe3zSWohYBQFTk
fjcq9+SRbqrR54m6mAa76Z96+zGvWBKI+4+zf1je96c6sa6jCS2QV+eJZORisfkCd44fmnJBghHq
L1S5zl0nsnDua7Ol1q3kCbiCC3B8lJqeTzmpxBphCDsg9XdoJfzf7eFG0Yu/XuQu2/nXe4h8LC9F
Ylkyl9rB9lCAhqXMqFYF7RqXt1bhlSKXRvUBWi68juLhUdxGfhhxKWTZAYeSXJ84Lkuq27ahm5j0
PEFFGK7Bq8pkvj6u8oV4Sz1MOLGjItm24BXEJeozOKMQl7W4OV6ZubAxlPsFDrqJ0/MKMfsMjpfF
4AAwuG3vMpSHwzfxJ6RXxxLjBanwf6OAKPzjiibRH7ErqpWBnwTpmJClomgdAgUcI4KCn4JB0xDQ
09in2cqeow0ZTXDZ+MbsbvaqUGP518Q+QDW9O4mIQvRPVPQnUOvQsX53k+hWE0ukZSI+0Yn/oT/H
0KzB9kH2BO7wEykyoQ8SW6zNo18QbqvTrEodI2eukE/SKo7bkNifpw0AMLmoow27W/DEsV4P4h7c
AsIZfcoIzY6vFggqU2ZgIz3DOaPC4I+VPnBO0Y0TuOQdRuwI4zT+3pGN5DtW/MJkMnaf7ts3Z/Ld
3Uk5a+FnlFgyF0qCwOFqKRKhmf8qoiZVMgwmfamABeBKOIEtZNu22nJ9xnpBU2FfbZDokFeu4BUt
YowWstUrz1LSRb1Rrw+6WCqpOkyAUV0wprny7LIvh61yG8u4+qyQcySYO6pZpgE8C/SoK5K1P07p
xSNDaQgStor0FWyGcORdX9ejATY9D2Mv9N/z8QaqwyWUOpOWaPXgVHvWeIzoIJ/CUCS3/qfxR7vi
zcoKjB01rfurJ7ocyf8JvEugkuxtk6ibY8J4BRnbcQOmHKyF/FT2WkTOqq576hGaCfASSfsiWkJx
wZZFu/Rv0oi+Z8SwGakuDLaI1YkNtzEW6b7qUjBCCMeosfa++WB9O+aMMu10cQ8K9wF3qsF/Dq16
+m7Mll3wxJwfQvWNuT3thyMpcJcc1ovFb5GOiNI+ciThoEVaj1DwOX8KCYsJZK5wuioeWnO8YcXs
fnSi3VApjo830lfO8+AD3xE4CWy7hawHSfEnCS5ie9haAAcBxQ4nbUFVKyU//fi82y/1jaDNM0m1
ifhbqeqMFHn/ReJNoXsO/Xv5WriEtaznU6iFdfX1DAAj6IwYjimA+2uZzyBoBWEj28NnTXyKpNIR
p2muqsC8JFz/0UeIQ4/p2jJer9efkdXuW4IXEJKAkdE37rTbVY79+xI3NCbnAN1/NGgRa0JOa4pG
5bVRlbbUpRTwLKbAklD3RnMP+rMpc+cvoZLqqGKH5i5QGI/V9kWTMXy7PcuZBWn3bRQQ7D5KMZ+S
h6OqVwGgwOhovw5yUoeu2eMq8L7VieImKhfe0LgtDTkihVep/B1+I2EqNzHFEulLzqLRaKDUWzE7
RMfTjk7IniRdsKJx3PbYUVqChLXvnvsP0QRAky55+kOwwbGmyXVwYDiberFf9EWGxX5LGl2YCuJl
8uuRn6xu7+c1K5eHIsBN8gn0fMLO8HRgJFg/UEb2BcjWhI3ADX8An84CbQDP4oEFW2j7cKH8R2wr
vs6xu1Zfg7z+sv5dzx/pPVlKjM/QcZhCdY+i6zRLFEIqqJ7SheFk4omWuAuRnDTwNKNrvMsBpV7G
jat9skeaH8NDVi+F7lM1zOL+XVqDGr4sX1GMn3eXevrAGGuv8t5su/+rQEKz1jZq132qhukgs3WD
2VfVDDGrIzJkXYXFxSaO8sU+GZTeRefMs5PF5HbMvyRxtAkVOI6r1BspRvFmEAhly4Ko3aY9bG6w
lCtYH9XEOSJ4E7A9Zak0eRfmZperc04l2MhT/y7/XkKL9wTFbcZ6SyoxlW0+Som0Ztp1PigCB9Bv
5eSFLSQQSWA4lub/CSdLnHv4+WNw4aEt3jyr8kYVY9kZXvVyFXbiv9E/1PjSl54LTR/JdWrpf9Dp
vEoyjdq6rvchpyrSApSUYnGKaqaLFFq/VNKsSZMJSdo7A1HgenkbMt9iFrhQ+wVe0dsjhMrwaOLx
uRI+zk1S2b+XY1xT3x1iLuRwbh0WFgslUtAbHoSeOGlnWHSiHge/hZtPtBTsbNf5+IV2zqxI2ex4
8yJsbJW3CfRB+/DBKmg4oQh6nX/jruO3HQUtycN98su+e08LAZ3+8MnpGiM+HLVuTmA74FiVDvjl
qjPo8BGfW9rCcAtB1nspP1OpUUl4C9r3zpuF6QwXYSlGmE+RRPnfAiZEHroCKWT5BRaaP8AaQdKa
YXPX/TxLRT9G24XWg/R/vaVF0oFXnJhRH9wfR/i/KHtoo+H5XKzVxkUN6Qw2z+mN8Xl2TK7pR9qY
b9oPoFi/1ZgxFc3pj7IVDOsdInvPF6ovUQzd5qATaFJbdqFa407E72hzZC/njy85AwCvNPUIn2f6
RxmF+tZ3S+bLl5kZtgtcDvkwCB0Uh6I5Dv3Sv8v0+BC/eaefX/mkQaw6Rhz9W+x3F6XJ5yyBKDru
kaXEPq3iyQvcRGYVfGa8NrGVbOE+/vWeq7WBompfYZ1Jlf+6n6PxsGHwW//1AtMNY9uhA0QF2Qcf
pt136pjgHrkIT0na++jY/uFb1ArvY84+p3JXk1BFODa7++sEJgNGMGlUoSRsIuYxLsDRs40FmyiY
1B2VXnp9PSa5TF896Eg06XIOk1KaUlHQLkWb2KqlnMxrzYIhD2AD7svUC6xEyLs5g5GGimePLUyS
vgRBGOnYXDBNriWTryd+Ar0fivKALNVigpfJG+L0caq9a2I7D4bh8QukNLmniZtwD/Hw1HJ/JZE3
mABDa77nokbeeIA8+099jQ6OvaNR18u0iaeP3lljMtdPfeHnHx3DXYl4BaAS9/K3u4wXY+gd5Opm
wOwLEEa4bnd6fU0s6CkclNf8mVkloUWtiYBZWlbt87kz7TsjDgLNYHbkiIl+XBsyaXOXe2nNMM6w
6jpMQuPQTI7OfCR8UcHPkbc2GyfbzUNfhN6jGZSq09dans6xLK+2R8bpRUy6Jpw4Z52ZiHaAINuh
5wIM5RZmgAdxLNdIy9v5O2cO+t5bAM3oyzJy476caUQ+lU4QtInc5TvAEm5jIeuDSZKG67h8QYsr
Cqb9mFfRoG/jl4T+I9/AaUArRZsKRYjOziB1cVRO/lgwSznZkwA2JDyEPV44DdmSSFQFj4jt5oO+
VPwWSyJ0PBv5XNvZ3UCYuNtK9qL9y42UEaG4TbQcltToEZrka5JWpAeHPWwD/N3iM82VCDrU9MGP
IkJFKXCT/6P1r8JwW26IyoyoZhjFVJOqpjozJzPmugD9vHUqOJIRmqyhMxjaMXzOQoKsfX0PCYWo
F3No/OldNx+lNOA93UVfdZ1kb49Btg0bdShqZCF7yOfqR78jORCu298gaaftQcgWLiOyNPvna17W
m8UL+sbjSsgLIaIvd6qWjh8xkqyrT6jUATCgNVQoqClk9FW06UNAUh12gr/K4pDEqRVDxrqIgmAK
RSI0OGus3DnuIV1z5fUhRmj8w+KA0v2U2hvrygs/+JPkjIy/5cecqVXq7VoY+h19u8td7Z9FtZrm
2lR+4ZBzvOvDlbc3cnznNr/PH/m2iV6QhIa7ubwqYnGBH0QyOO3oK214s93xjgy1CiBVJdg8zmI0
cCGXEVXsrOpBj/mDyUEt0Ja1VK1KfA6azS5kZKjkq71XlmUKvJULbuDshu7Tgzv2aC0f08fJK4EI
LUgySV2pz16I8fqGd+/L3zhoZec0TJlnH3qN2midaL/dmeuVU4HlpO0cp3trDMvdjp0FZrvsw8EN
lOhOxCNiapJZhqEHfr53Gd59zrPttbBaNTd4BbQtrRHePLHvj6ArTX9Ko5lf9AK7BrKHql2C86pb
nUSKZ5IKHxmyps6LrwinQiOgFH2sUefjJgnh3ARK6HnM4kJKqQ5upl8zJO72/VPAWPz7XYSKovWa
Fpp/M0rBK9XuSaVRwa6dl1VgK2n4o0QTxS5J5RffD+5Zy9CpYAu8PsWoY6LJbSgzSE+EnZQYb4mp
lu8R0jkeMJryV5ocK0Z+9eNZgODF9p/Hos0YlKmGC+0fZVJf9hN5Q8qx5eD1MPZ+L61aSqAv/1/0
fAzb6E67Nxc9fc+5aEcg8903YRMJpAFPnlDLeAY25SRcV634qOkF+depF0OZzNXK7ww5ugmFDjoR
VT6ynOOpytTKJ21f+OCkEen7kf9lGttuXW5k84xABkmrraFO1PmTWyJ8ksOpqvk6OFF+EbT/Jhws
8GJNX2wwyCFDB3taYNIXx2Z2P9S90vEbTZpfuGA2GpOkrIm27+w3N+Vx8zrLyunINCJcCuxxCDi/
88KhqBZvD8YEbcicfM73ODW44vA7NGBfbtkVYIIbCzBse0A8d/yHV7KNMsEybB5CDi8eSVJuUjH4
tcC2doQ1OJTL3vTtNmTQqZuHaPhRPDYl0YLGat/BG3PXSca1sIUjzzEYfXOpgoiy4MXrHq4Gc0rQ
kkWjmv1im/agEKRQotXjD2Z+6nYRSPPKQaCUhbjznFeLoADwzu9+/RTV2sQPd3GWHljflyAKOaju
ouGSCnbQqUp79I/8dvRFpPH6qnrkyL/Z3fYAwUv9jpbwX29HpAO2MVXuSeJ+bON17Gc/AjD/1BYs
N4zC+qRvV2UP3a67PgCata3WDTUUoGS+Qib7hsGslKLg2LJAZf8Fnr59TCgukMIiqpRwm+YxKKwu
X5o5KOSyanlLTE3ZO3YQ34b4eiGlEpGUhfldgX8o4cHeWa3PrpC5Qb8MlNULLTyej3WGOcamsSnF
4kEEuFxAVeHyBsu6b6yV8z2crf8FOknmXk13P+5xIRUt6tzWKhMhA+ieXX/k3podNUKwtUARxtlu
FHs8cyp1o5DK9RuFTxooNLfFT8o11eJ87YedlL+JAev440O7wfqpNt7vXTYtGBBa4ZPmKKayj70e
wc1PBEZWRF5zt6yzmBtkBR+y0N8ETIe/Vrefrwrvv5qEGoKW0SBsXqViAlPU7r44DR92zJjoVUK9
4eKwIu70solEtoQONiv3zkEV2NJt4dEzMnCVK6wyEk+M7YEiTO6ZfDj+lBo0tUZWeM9/hLjB1cEL
KPNUweAqSd/Tm7vPCB5KSy3+6DHvWhGzgoqcN24Ge8/ffXD/h3vw6S4nopmwINJq0glZueq4Ps5m
Z5tQGeJH+jhQ0i/ZjWiHjLTj5SEiEVW6fr2ZioyMLzF4Elo3Aw+kjbfE1jex3B/JZmP7tLyDwr18
D0p2GBxJjfxU0ZZ69rMLv+7Sr5uH6rb48UG1sSFJGOuQPGnZtUzLe5ZR1qeCNlJPLtNlnazg3TTZ
XI7bmNf74Ks0czH5f2rVyhkQFnNOUmT1HPcFUykq84QuTN64KO6yB9CUhKNikmD2JG5qwDtakt9x
aXzgI/f3Ms8+5LWFoeyBhmDOxnFdEocKDmgopvcElrnmth2ClDoDsdec7Vs+2Xrhng5dP3GWgazK
TXauQhwpALp4NMP+cVLIYmH4T/W4jVxlFar4BpKUiBCm3v0YSwuFIy6kIVfow8Pn4/3R2g7MHs+O
G3PWCROaMX2J93tpH4kky+ibfNlZD2KRhB4Wlsi3akWOo8gGPAjSeBzvWoIBsyRdVN6hTRh5QK9H
PHezO5hFYGhEK81rbofwU0jJ0O0Kx4eoGSadU7c393HLKCGl5SLK+UybXz00qkg9bHOJIZPGNUoR
QUktqiZzdWXvKQ7foP/qAjeH/ZCmMh+bZzbMVyLqJztkI+e/BrPRueeLzkk0+KfPwnWok5xCCZR2
peBWciuGi3Jh/fgJnkRZUSGFZb+xDdi1vdaopIS0cNXkqKChuzRrywqgQX96tvdkGSwwDvyNQTEN
imUN0iVi1rki2X1XacSN8iJSS75xU40ls96+6yAJnKLsft6VVQpWqJZo+MC3ea9hK9P9Z5XW1YnH
n9ZFHQmkrM6XGthYdgqmo2vm2wzGH+/4BPKpZWd3lEVRhGQPCxkxlXbucyirSHdIWXPukCfm4ypk
77DH4VEHlSxGo/ZvYsLzTkB6hZNEjGtlGNgFhCQlCQn1LBe00X6pZv11SJluFc1YS+gAdCuLrhoO
TKzd+6jfWPq+RlzUqgXrj7OZhnzi8W1yNr6hSJPOmuHNzOsa5g/HZh+u/Tohss3P3oqpbCI9VzRl
q64so0jA93dNHZJd0rLJetOmyStNFlLhswC5YoZzs3UGzBrEyAbWFcq45Ypsnizy1cj78Qysri50
m8Lhgic7b2n4vvlBaYqxNHQm+VftkymE1uaUZIMOHjGJXCfW3YiuAJtwXtUeVp1KcEie9BWIKQda
tRYjvq/Ve2lX5//ufppAw9zOw8jDIm/EIIMOJ0WVAeUgVMsWjDJBhZOo0CvidQ7QpztQmZkRD37d
CsvlnOvMQoKXt0r04PhdI57hfPnijMM9MKJNaI1E8Kh8vhMA4oK4wX/7OX6Aq71yP/2o/cjxMA5y
Kt2qfTkPd+HnSC/wRXBKT1j9zq7Jh3iT7nTWaOlodwE+0YKFBwKcRaPZxo5gyBcRLrPHVckVrLfn
sf9vhzunOJkvGWs2NjOntkIuwoWijFZAd+c6fMyCI/hIfTs4kDmadwcTaMH+2+wnBT7PfZX89M6W
9H14/DrjMKazpy+hpiHR0UXp9APEaaXjI+K9YKPAc/okRk6WwMxor54UCGDjSdCS3M1dGCOkqJkZ
UpoiRTvK0UHWoI7qECqElTtFqZ935fWTZfaz1jDK6PAzmnizp31bNMszOqQ+SgwLbgIM2NZ6kL8+
lXeYptqE3BK4EuKy5Y7B4QSxiQO/ftrmkLjkkvyZVdxnm/w2IXX6u7b7YW2pQfd1xWBX9UcJvev0
mfH+JGLKJDAsBaIW8J+zqHY6klUL2El7RCoZj/a6LDrOzA9/7cVlgtUSwVgUWVzjymmFkm+YJxGU
S+cLr4aknPQU9XB1fme+gb0zVR87HU8YxeK3Q6ukFKCn9R/U16vpkC9U/l/HgvnS2TdE0wxqvNJW
LgBDno1kjrSzanj6oYGq+S3u9q8hMpClJFKebE3CIQIpcAxW5iL8z0q6ZtEC8b4D+HmdU0fyFilA
hUtor/0bzn24NiniNpK4+d+3/d6CiXdwqi8F0jCQJT8hHW9u4HKAfj9MkN6zydJv3AQj6ziFNZ5f
lOCEd0PaeN3HD9adgreO2dxYTpcdJbFcDrRv9DPhb1PEQlIP4xm4LZzALFFEoJ7vdkE7BnYNhHRy
D+JT/WyAYLsqNudNkbzQvijtWOGc+ngm+jTSjU4qWxOg81dSFHj2TW8Wyt9B5Falm7wfUpcX90/S
0SUVGi50nvLcIl9MQLNmqHPhLzKxpCHrFX9pROu59ZwvebfZFy3kE7WMNXDSbgLTLMsHMIW+P7rs
vHA63JhztU1+NNCG8pywrDsdswydxLMZTXxYWVjzqPL8jTod9qkOaP/RZYk0S6PdNDMPVnt1mE1Y
8XPnKrNnbBSxHyI32+SshYxrfKobId2tqoZyM4wQ8CMvAsD8VLtzizPCZW0gwniTZwInW4YFkaMn
aied9S7sEfD9iDiix/WZM1GHJ24B1zhIPWuUk+dZSpxy1IarLSu6462PdodoNeWkHDuL1nwLCfOs
sAcs8Y589w2fUNQlmmk/mi2TcghXsNiHUPT7iZiC+T3KKretQdIxsQH7H12GILIfcKkHGsNv9Op1
7iTGb86yTzpM/2WsuPLmb3r48nbeForTYzPE08ImMW/wUYisV2Gn7MwQ3usI4peseL1LI4BCVEkI
d1HfWGBsFYh9onnuXsY//ti5dwWhR0aVjlL08FFlWF/Jqoe181p0LCIHaz8/zSvE5PtiRblUBzgv
eG1awaDnpl/oNv/q+BELyq71Vm9dHt+P5P38y+GYqyUGhSo4MKJb8JQDVFYx3Yu1+wK+VCQ0e3Tn
r6PgXTQQ7kr/N/0k29Af8rf462KMx26TA69R/+qW+XBdh6bTo53GeC8kDtc5WBpdHJwUuKqpXL9Q
hiDolmJZIoBhherQSTjXsa9yjM+8jlVuwR78oT7Ktxi107Yu/s2m1sLbnsMVcGoiDMT3WBP/7dxW
JKlf2qeqZtp17IGEZe71huJLj4ogYaU6KuEwScDyBheJLKq03E2kFYNbptF9x5wZUZR3lxIDKncS
310OWGaEgTUuuAlPa/8SxEPPtGkSriO3m6QKwV3rGyLrk/Xe3v56VjFwJVNp7RyfNnaGFpWq7qUU
OFa+5iLSCne3x7Pmsxx4x0xXskclXbPaOnv4+iCryoW2ivpYoOjQRRxf0HIuiARKIFCeBa1UofcC
GO3bRKb8IxxHSyJQ8yFavcPQc+slTQxkVpW8NE4Y9xRjlAtsiHvXutHWZdWKNPrvgNCKp8vUE1QC
30ZQCVXaIgC3FuYPjHODlOhyFbV+Pvzgy+X2RAYDFxbHWnUcXu8vC94MYjCFfndnVvtGwk5s5U0D
hVJiWOmWh9SR3uziFbXXY/Opd/jJpUc2kSXju/NmhcKmIm3lUkf4lGsXz7tJoit/fHCXn6gdGk8e
An4yB/ExFWfFCBKjtZa6+DRqcsmf62orxWG/2A2IbD/ybx2n/Qjc5ZtfSjoSo7HwtB6wSy7/iHGG
NXA/LzFbVBVFc7nU1j0pT1Shz55kBg0zqujSH1rCdOBxZq4X0fZpL5YU9gDmyWqUls2FrnSRnHdU
PHorkjES2Aznu8rWbGOza77GAfCRYZW8zhtgUByBu6TQLkhwYOpnG63tepMdPAZqkM1Qmt4Boh+U
CJYKPI5N/e5XlX0bR3866VNwNd/zIO1JHyQnuImrbG1r40eizzPgTy8sHEgj3KmeOp15lcMHhJtA
A23tQVFDda4LaGIHQxhiauxWq5agDxvOncgwFpWg39nrMq/w9H4v6iTccsUDDgeRmdFYKrQOV6/Z
EZpGs62aycoNPmXXotdpz16jTVSMi099ielVnBQFgKP6ZwkpUjUyPA5mZUAdcd80hHvkVmLa+ciU
6+kMxYoCOwOIP/815YZpBIDuBIrGueb+/M1pqpwtc6ixpidBIAwscWZNESN5Rmnch8J7BjJzYqmZ
I8cZFvk7AdXhnG/HlttXqNrJalM929ogth38bCEGiY28REVopF08mG0mr5kUM4GSQ23CGOJkD39y
PpyA2o68vrH+9TbbSzgwreI/zSUe/kY8aeGevwEjO0ggaQq68T3Hgj4AJoUqbx844I3wlCL6ELft
YlvVKs9wiKv8B4Z34BpeavBw8f6viUwoEhr7Qd7ztIGz5huHPJKoq+nwg50WuSYK7zVm3/tzb/zA
yzFuwulWHfK2FRff/Ys0WU4KTb9bsTuZMfj9biUamQYqXoquUjsoghHmrf2NOkiObi3P0zDVS+UE
VjyRvT+3SUcbOXR0F20njCJqhxWBzsHPuiiXGSMEBKvXFVuMsRsX6YOFaCrjJ+OY/Yk9lCAZzgSg
xyqCpVpsDJakescUMsKSnPEm8hyH/DDbzb8bpLqJMvl0PDqnjsw5sr00x+s0z+4l03lxoCisXyN8
ZCVAQBJ6GjIHTP3oYEORiZuRbETLowZXQuVlcpYALkpmrafqm8N0xvYGNtU3KgVdX951td1EFPni
eHYazZNIfpmtFcgPFdmauKMh/9UL0yrrHPQmHu/pKVX0B7YunK0nwUvbo0J5+amzwVHRmwMda0QR
gnL0QI/yzhO6TsVoql+ND3St/lOKMFFGIXvoQfw72P9N9h/Re0hXKtjUX0+CDoJo//5M75VT4hHg
B0HBGcHANsTl8c2yRJWYYwV57gSyLnsny/YILvRh4j4VfcgTeB/+XD3gmgu6hlzmiMvdi0AmwsDB
uZ8QJ9dc+fX1QOOMZJDXDaNE8xJG9+7beHXVRG5SMaMN5xnhAVeZHtcIsIgMa517sgiCRdXpa38p
jjTzQskF/KaoG04ct0u8x7aGDgoCf4nbEygG9AzydpD4kkHG9NEKx/oM5N2NlzqdDTR3vMajj6Gn
VngCCsGTNJkZjlk/XLY05c8len+KrUjj4cVgt31BAcBI82joprZFqiG0hxXhfoBVENH6B+EPtZtI
M+3fGCJRUGjh4nCWj0wfEgqz95qrHZy4qjQum7DAGNajDxCtN0jKnXJ3U5OkSukqLcviagOCTfrR
sK+NnpRIBfGYv2YENQKa1HVcBXQuQi2ZtGmh9lX0/vanGJhyqaW9+SE7jBhdXkVry7qQiOX12SzD
uA+/Pl09b5iOziUZXoZo+T9ZcPcLYi9CzG2PQv6ggMpIyQK44PjG1JkknhqrqPQKlSiBhmNJEC7p
s7w1o9oXbUKaiEUymrEg4wz5E7DAJRIVeA8iVImVMdNjgUGW4H4tWi/YqDEeNoWOvWlyRV+vT7eY
RRkgnUuxyX+Fpfdsadyap89YyBIztlISSVx0i2N8WIyDvRx4JFYZkozhWdXT6y1HF/SZWmPadE9a
usTGpphfkTdOKGQIbyxCTfnVhCbhsuNrVGF6cYFGwW8osKMO/F+V0TIm9BVyFXpXVjcS1HyX9dAQ
0q9zAqcjKP1tOfG3KCF2PDa1wVlgpGMfH16cyZo/WU5czkbXDH1FPRMNxdP5Tzd490qRvFxZB6I4
lgn33/t04oVenvE7J3XlR4LrywqBOVvtpaDBxPtuLDXNX7sN+qaM6oPfoHruSHVGGIplMg5cLON3
d3dkKDp9ae7RurjDcT3F59iSGCJXPQF5TUtP9XKZN0qtl5cmLkZVzFgHj4/f178kbyNUCbXjQsml
EalBuqhzkHfdb8pkOF2gq+kcG9wps0/XY+cd8O9oi+2gR/HkYd7c/vBMNCII9Mk1NGU6k1dSwJpc
CaxAtVUnssTCah2N7JVRSnYIVcnyrHSDJQeDkDeIu2IGAgB2jQqGqhSjCxRqo8V34KMJm5/5irZO
dSz8kS5veu2pTjWIodIy/c39r+Kfk1uJrr7YJ8nTVxkcxUbaOUtnL60/HxVSjGcLmcT9ntozkOac
MZme1Hi1igfvaOoA0WFPi7nNHPTKPgBcvwykjvesDlplkRkyhUoIi9u1YCPuNZrxXRpAHAEkB53y
ETjk2ym7J4gQKUmUnmPcgcKa+7TIVnHyGI8w1Vv4ooRII8eSIB9+Dq5WgF/oL+oXeEWNjbPDZywE
QEze7UYPYoH7RIm34gvvUnUbfYn5T+oAWWJwhX4sg1jUU3fy6c/HqUGr4XVF0Rt7l4fbD6f95RLJ
/QOKa/7lb1jldcL5hlnbsq8h/eJc7RiK+3I0UoWMiLSiKnbexsuViQb1vuvZBqjgHIb9D983FW0U
ji5fHTn5Byn/6X31o5GA/dJUtp18WOxA6r+nZEOIjORzNbCr2J55OFsRttZmaAZro02sTW9hZIZo
miZWnPxsI+Rh5xOTTdHXgzlznX1Jav9GTMViG+o81pTGA7Yyo+1Sc8TfK8KSHEQYyeSS3+SYNFyU
D/14dY3fLVFLKcyoyvkSgzz4NTo19ymKuNspV6DDW8bPTmxU4S3HMJidpBg4vt6L07F0mrFT8pTc
dZnJDth/CadFQBvQYpDSBJELeAzDECtfC5sckqoHAsZBbnfsmNkBMA40jV+ksBZTFAi2CNvWc3F2
v1Xkohzoo23TUnakFop+kf+J9gWCG7WPn2tLu/cGDxZn7eeynUboZjfGzvjNRg7mQJ4dpnNw7mh5
Fvr8hkseH7WgEQmNc0pBQBEw1FySOK2++7RUlcDvVDyNegU9SnBJR2rebfhXqrtD6/CnYb1B2jKN
j92NYgXBGicB/xXCsFtduIITe5GMvNrvaxZ8tIxFDck4xvUybzVhUyPFHvhBggGEL5gq9ToQDg1V
B11qvH1Ey2B8vV06MJM2uwNxyOwBnuujT4I3pb4Y5YviVzxMF5+LUbUODOv8A1tBaNeKIgswk4+x
dqHb9mPWsnR3ry0sVlvL6kMIpBhJDfunpaCFfH2hw/BL/lT26Bi4dvqut5+8PnEF6GLJB7pez/IY
UiRr2t0CQ/BcK4esqBEImieAmUqFuRJXVYafRYgdOfPub1MvIEuayFZ4nkQVzfSkPMgaqpLaJqQY
DvUjTU7xpugiNTAQRAlug4ifJmW2MI3I59t8n9/3vz3iBzzAfaSp1WhwpsP+46k0wVicgl3Q4nAd
smnq/soNuwSw+qzBBjtFFixdC9yOAz0u4i9xIFXDSSldwnZN3Zu1uOi1JFiOVpH+1Y4n6GQGQhcS
hoENEQ3l1TU8YjpnKaV6b49GGh86X9LFE+kF1eR7EYugUA66UXFUEnEUhZaDBDLplDhUVUUwoQD0
DeNtz5W324ehcQPPENDZjlSz5jkMmRjgbft2+tgf+lNRM2Xg38lyINKJqW5S/AqZFE1azqyuIGjv
5grUqinf9xJIUfJHo/aOcb3Z/Kond3KIegrhoATebPuCCua2pqNwvHQpXr8fSG5ubGynfArC1CIC
36alqHp5Nvk0vy7FDVsA2yN8RSiEFXJ+YpfBkVTcYOI226ZlsVpaCI3GmfkOwltui3OG8S5/KAhJ
zpqqFFFOADSIpNWnl9MGtxDL0a9irib5XNfU2ZHB4+AAEO4DxyyqcXTWGry4o4yU2ZzZxSnHQy7Q
UF7TzUiesRPXXSz0/h+cbqSSkdNIrs5qBCwcIxL6pHgc07Qo445D2DVwIdE800FE53196FZPSwq9
h8GqLXSviRI6GckwvspecZZ2mUcF9Aq+OdA4d45Q2WX+W/jnTHCIwC3eVudL/ty7hc506C0k2uKw
q7h2DkWzxEFBSxfXYySUn9vrMmq4iTqEp1BMtpOM9MUbX9qRjUwTCtOLQAPUtEW3A435aLt8PiQQ
aZ+rNJs3gqBkxApwh9nl0cLnW4p33Yz0IX2mlGk2mMoSnVD64f9NdMZs2+v6ioJaSC62qIlKTjlO
StpdGp4UXG2deTBPBmAMfDZfhlJHxbxsqVG7Gvgg3dwXzz01AtHER/J7kSHpljlzrf+0iTKXTmpL
k1/ninD6Ax5DuQv8AvSd7/bpras5PCvYjyOyA/GSOlw+B0P0svDh/xoz3iY+cSTdsOtJlS2QoF5Q
5GM+YjKcAEiDZA2XYRm7n7A9BfPDEiHCuOijZgWEQBgO4nZXopXlaYTrzJYSNWSJO5mqudPOdwpX
Km3f4QHbT2sHT6TuLqQl6moX5NUja/ZXSXnODJJPULUXnsyLVX8Ycw+AQggDQud1KIPDcrhZ9851
KyWAL60nzR+207qH+ZwpqGpvx1UbDamjUL53rh7XZG+y4trwRgw4Cb8xionx6GtFJn3uX+nAjHTL
LredbUANeO8Tg0m8BdekRdTcdLv6V6tn3p+LAkg6yUi7UF7R+dFskoGJKWO98p/c+jbYUjqXNqI/
8Rd8wwVSjcmv4jSBH5oQn0puV2tjAvnjfBG2ntKo0F0cxlrk65lzMkmTKm8Txhm7E3/NQzWbJnSq
I4ffAfOEuG2Jian1UH5fZZnkqjIygnyd1UuaKyak1sYZqMfTX0jgjSNs1Yg4DSWtigkNorrnHmKM
3ZZMquhNCWcV7Hll1RbIHIzkbqi8hi1xlPRlaGRUjOXAMMym2OzIhVCcGfXu2aQWk5sw4friOKZl
1pXTYw+JjozG/5lmjygPmfcwsx+tC8ZK3BGmsdyS6Lbnz3lXEy08Tv47hp+HFKnoF9KmQa4Bktum
66yf/MWobWGmm+EoqaLCRg7DRi5gqaNgyaixxAmk6BZcGvghGsou44V80KDxOvDodlBxjE+44Xmk
gGADeFaZL0nElEWJUqjOTozaUu0Lfvs4+ZN0wsz2LP/lr2sA/tSUzWiU9cjGAmb/VkS8HuNUty6Z
cfpI/GRaQlKQj1BGRBVM6u8NvbC6JbdL7fpDAtuSN8APzeVDRrS1IGELArPpV2Ry7/P9rJlJECz1
sIpTdhxWxR0pgMQT11H1TgdZizKeGEleaQzEoTkj6eFPNH312V7QpZr/hUaU22aAAUtaPypqJ1iN
an74UWwlworxT9eHvVR6unt2FteYP0aZZIbRiCC0jD9HRnpYllmd4zGTa9BoamQBOXeaQLuwB8V0
AtHTPLToI/9L2JLYmOmUxyyZV8g1FaRK8HANLwj6WXeB1hjxIY3hPQ6RN7vQc2uIFtIPcKT6TULc
vRpRl75lKn+y5TlaZWsfRQteWTKxp/hcISkcqVehfWBf6sRcDXre5RXzTwa2DpHm/+RVdOZUkms3
Vn2B/VUWpEn46BjDKNBnDi/jv0FAI23xvAhuB0CA+9ajaE93fDTWrxZwa7DiUUB9lhd26shkOlM0
i/Q+PET/DGcVEciaubXnTTEIPidq3T99f9tPPKsb6QKANkEIejasHvIqQAnRUOGK3Gq6SC4jqjRf
nvCJRYYfckiBrmWk6+u+o64QKdF+GpOk85PyjbkleA23yx3oC5GL/QxHQV0RDD2nFnXUdVP9BU7j
Ns/ViOuSkEd+91x2heGnqduToao20lxA9fQEQuDtXsS7fX7C7zMgN8yTmB1iIi5r/TpVcz5OdX5P
6954mcO99Wj6IFS/ngfLo85UhXMeqaEB6J7XgvbJAQUIVsouSOx1ZMMGCDpZirhyYCIBwLRrVgbX
Nr5AHSE04RugRyz90nI+MgZ0FJcaiMMbngtu+Agq9gOQRfPKuBKVoEVujN6pKFknxIQrQ4N8jgzc
js1aAKGelEdqa2s+prYAz7JyIcnC57iq6ONVBgrC3KPbMRQhHrrrUWXqaKi1pXNBmN50FJMrH73i
yfXXAZAaHNlCKmvPqarEuboJ0uWm8Xi7ePsW7dhVNt0M9/2zsmU5fJmnzIbMHouHl7YfAoaQCYNK
Fwoa6XEuXbEjoccQiW6PqM6YmZ7/vZStWBw2D4GIiNUzigRq7zzfRZj9w+rke+GbE46hmTDvqu8b
mGhjXr5s7iXLY2p/Pcz28+nysz42ObS1qDp3I61biPcVMGXkYir9ftjW1q0Xc5Qlc1YLQP0BUTTL
vCb8GV8t0ePtyeVancjaBcIzufjvyG2ic72v5NoRZM7VdWOmPPPsqmBZCQIm5nsvTZgZWqg16WC2
FsPeYR5kN6jMVQmHsVSj0Wxb5gLLINhs8C9Kizpdc4UDYvClE3JjLj7+nyTFJ0EZQPkQIbWJQ8It
t9HkM7rEqtcpxE9rd3Ws9ZjTlAJDJk131FZynf+Q9b2U25SmHm0/s26Sn5Wq0xM44Qjr1yoRaXdU
m16mdsYS1kbfsxGcthMsT3ma/h9thD8hJGPxxToizVkFyZJ4tj5Jw9JtQd2Aav2YBY/g9IhwRXsv
g6iU2e/vB+8dFE2LvvDPEI4CR/VRB7xinFFW3QcBRxWsxzFVAMBkLQgbd+cuPK5ZvC/v8qkWWOlh
somEeY77NOCKRS4fF2BoFGiVPq6zXXdmYDge6Rz+vdWM1Ld3fG8u5G9wgM9//zJliM8QM2NzqUAS
/GCqFbEwie5tEKrFEFgpWRPoLjCMnGLtlr1LSAZ0MSs/kpKU8ljqwWS9JvaEgRLfkxU1TH/RZck4
x+RABf/KvLKSbNsWm7ht0Iz9uizi+55jhwM0Lg16nGgpwTUlspgKaCitrtAnfZspcmpqziQJCylX
IFYDHGmUtB6HgRIlwH+i8VjPCUtki5n58+1IgIZ5kIFSLXJWB6KqElZ34oDSL6CS/6qrcecWqa+V
+mQRT6CIlJKWxCO0U6Yg4U1w1RkK+7nohGstldhD/OT4NRl/y79qoi/0fudvprPAY19hWIsXOOag
/aB2fV02zrZukZ1RegfOqq9KyhS3Y1TTNscoYXR3+aM2hxPDcvCvkOh/6kmQgXghDrifOD9vvQWX
mYnteCu/iYV3JkDz0W5Gwl4Du8y3uVvOAFY0W27lY1kOEQpdgIKlCc6FbpYpjY+quaHWwKlv9SVM
k97rwOwECJ318sPrQhsrnqoQo5ZL5urL6CUXJcX2rOoMcOQmXVnDlT5KcsOKlAnJYNS0w+PGuEDp
Ahvz0K8l1l7JGAMxA5lDimF7s4MowxaaGXC+uNP4iY4GW6xHWG/sulXwaxQPK8tShx0SlPmmEGJB
vFFV+2BDA2iQZAYYU+ujDpB4lAo1fblDVqdzMckHkbPHmPCt4HgbYMO/8iX6q3liseD6d/NrIyio
jy1KMG59+RekuQYlmNuXo99OupTI6nPZMFgyd2SKgmxs6phJ9jMcy5EPTyF387h1wwlI7Gs9+hX2
oUaSJtZmTrCSedzBxNWHUPhqlbYTuQyiaoZL9/JvMVk6rgpM0kPat2TmWopw+8klO7mtCJiYGTqD
nbh+NIGlerRbUVZ6cP2RE0u0d8NxpEoTKs56h3QTW3QySlmUwBuUezg9yOOOpDab0rnAHPLoxVoh
VtCciKSq1weFVsa+/AkxdRIx8GMEsdmg0YdiZ5seWo8Tvccnxuy+WAN/QgTYEEzc3Y4tFeibk7jo
NVvoxNq+/FtVI/x6IOnDXE8kv2KDkikTvwBu3dFAav/qA7c9/vEKG6nHePJ54/NatJWAajFi/Wa4
Zbu64Hkas74VCcSW3ppai4ZwxylTYHrkOTsNyAFJkMZ12Gk5zrf752HvD2aP6IJYWo+DBWYbbyor
ZEjh9NMVOUzMpCUo3cW6mZn6kJelYf8O/DBtsO7sxFxJkvxpLCSnIjg0PciNCGUs+Qrc73gPhT9j
/cTHJA8jSR39S7r9djD7XUuShdg5gdQW5afRWfOwm6gm4lkqjA5+OzYu7OqBm6Ni0cnBIe3flHrk
LeyrfHvABE5Ho9whLB8NLyEPMUG3CcQjFvnfUzxv9tH07nMetJIenti1rl96TjDikoo92+6tgqgj
TuSNog6JL/zhYJJI7SLNAR8rs01zsYJLZeSf8aBj1pRwmaTsvWc6C5YBSCikLX+Oqa3NvszwOvZi
gl+hdSvRjJnJUC+hRl5XK5ryoQLE/jaGCzxpKQeNrZpgKxYvNc2zaULY8qHg5iuAAa3QrAU5Ejjf
AF7O72jP1ezsxFF/kb4BKKI/VzDPkCRR90VBIyNoMiVzeZ0vfoAJeyOa0UFvq5kONrrK2PsQPaAX
DaWwUBgEkdNuADxQMxtoZmgvgRNWLey3uW1GLDJ+xCPtQs7S0Z1+cygLKqoRLprIzV4XX+R6dU3Q
4RnSPpHa/9lshmVhSl7iS05pf5F2rjtrFXL5e4bZdkoDcYopyhqiE6anbxi4wrHN50uqzxcxcUnf
VXw1eN1Evn4x5gTAi0fYoK9WuczQl1q1BCsCEUZEnOOHV3yD4PDw1pfszNaLqZb/LAJwKMWKRDze
ZeRFXMqU51N494KG38KVfl4JSB0WOhAOjefEeVAkngO8neTc7IvAQLiXqIAHbLu+Cq7LPkMJm2Hu
5+XEV2OiuRIc/B9Tev5UDjkSN8R3t7IPMZ5TbvTyFx/b0114okndL2iclvvtAntnNLcwMoIxUhMJ
985Shdb8BC3yAz6TJAyu14Y4jF9MOA3Pd3grCOS1EgBCVV7nvTFL8pnYKrbLVl3LMSSAAsZ/ObVy
FN+IrIV3qlZdJEc3v+ENiHHrjF3En3s3gKfdC++fvnltyJP5DdI6uQo3Cqrxuq94wXocGVSatQa+
S8jgQ5s7VWbntr9K8fjU5yW2ZIouyFh6VbKNSMMtq362+XRWyzZ+n0fAzj4SENbIZtRzdCrm2eCc
zsLzKX3N0U/Ilg+I8gM9Al8m5CCI/LCC+9HevgoI6VpjhtKTsTQAOBDsCMjmArr9aWHtUlGV+P2n
8qdgIFvLfvNWW1z7ovl9zAmHh/PNR9c0Cp7hSCLEqD3T0XqMC1nhSe0C9Pi/zUPubynb7U9jxxp7
a93BwxI8G8wuXxUyrh8fuq2l1gUWdt4EqDmmgqbNgChwQvHFe9mNwBGJFC/Sm9UdKQ6NQyxyEeSw
A3FWojJHauND+ShDuJhdW1UO5gNnodgkeU0ZraHR7BSlN/WCriDDML6iG48whBfCGSgb+fE7LP2s
OuA2E77jbuaxJ3b92Uq2wgQO2ICy53YLdUOluvDNHE2xIAd2yFNbOUNiSXa89EJGcfTR5wrjie7K
V91jLeE/axtZLR8VAU0gFP1qE1OgdSYJbIcZwsZJHI4xzhO2M0B7tMNthzMQ3RHmUSnDBL57fSjJ
NZgvRT+6n33wRldp2nfKjEvBffv+RHiI48n9ILRnUT3h4jocjdmmijrbPPly4J4Cgo4WIIodpJlH
kSdYw45SazcdPj+bnUh8LSwEMQywTPVNP6lgiaUJx7OtmntJ2riuepSEhg4WOAkk+csF2r+nyBbX
IDQJIpJs3gaEKqO8I42fOoUi2vsFeRwvdXqUXLC3y4vGFeymNiDD6iyUywzkNZXl+lJtMwWigz26
5Xlig4AnsWr34ivziG1DZMqeYjzdmgJK0uOlWdbiZi8Zyr+S20cxZ2MSq8ywtRU80MAVMjbNkrPr
1kAHFiVQ+IF2TS/itOyB16VoCc1vQuVzGn8/DjJZ0or1Nqi6TLABLCFdBNzvftxcHgB1Q/vu8lzV
EcXrIOUxpN2BTjfNer5tOgHrzN6us7tRZwDW2Whsb7tRc3v3fACV4ynh7TpWMyOVzfXTY7IBv/kI
CoIfGwnYRTVHWOIJjMVmaaIs5Gq/lrTBfOWEr5rLImTZ1IDbgw5nd0jv58DrkRgID104+VPrKGzb
u6gybJgF6zeGREJjAVt6tMJAJVzsdoX3c4OxGOfVUS1a9R6YXEuBtaJLiXPycU03tIHqzMq3p80C
TT3kQ56r13veA/papHpZD6XAsQD8yeXwWHgYghEQZAuAAHyraxK6Ewhi2b68K9LU2nJap13xfRTR
9O3G9irTZf5wjmQD+8hK1yYpdLTw9Z8hRLGrdH6jSw2VD7oK1ZqAF/mlnhDWs7Ej+zAhET1x83Ib
BGCdk6aAtaWheuEuqCVYLHm12uRmntF81UsTYrBApf3VHUArupRnPUdos6U5mqpTHqRm6FKNTo74
v4O9zFW42luc5oprbSkYH7+dBWCS3SrhLwLr0YPlmMx/iqI4vf+JtpYRXc5U0yRhBKJZskVmb2mX
lXKzd4+ExMSvS3Elb0UmTg1PUVjeAWm+QDvTCBQY1nDtrq0GGk4GrfIhyUcXV5++iWV5DfsuDNOi
ZR9SvKxsosR2kI95BNzN5OkWkEApp5sZR4CxIhGpuk1BJyXhtlI8r+YKkH38MxeyvCtce3qlti7j
N3feAppDlbiF6644ZLDKh7WIttVsLrxTPVHr5+MX+qYrR4j/vN2+BxqmY+IDdQSsaO6uDWIKe2vF
xp35eVlhcn+bSEqNtped+fYUUrzJswgofFboDaGHg0LgioF4uw7GCfOniDwWy9d6Hrelb0v08zBT
JQK3QPAN5mlPju2y3rwWsoc37DO1N71qPO2RCc1K5ZO8vcJ3BCDbrcA+T03aJlXNqmtJM2HK/psO
TuKQsIKEKICphzLsq1OjdSy1t+xVResy5/gJxTgXqWi42FPyxb1dZOW5F8XRC/vYjukRm+Greuny
XDgqGwA+T2iKZnAAEj1gGwDN1fU/fptK8pFiHtd3J93Rhs1DCM/T6AtkKHC6DiHVLsgj3dIRhoH9
kRG/5OURXWkUhhtQ8L0a2Dgjh7g6uYXKTTiTEynP7Fn01Xl2rUFfsF7BN4D+N2m0VEilFgeneItC
afK1d+9ZWnaZ2ouHevePk0gCTMx0rzsdlP49BINf2LzJXWSrf+JAvsey6r99aAKj24Hb4w5ZHzid
aNQ6sb1Yy3tVA3GY5yDTnEycOtY5pxyu1b1eKVB/8evIMS48FE2df6tCBWgDEZ691TGzt+UkMrU3
IRVdv7u7zm7UWHc8i0TP22tecnesAwtmn4Mb9TxPvlQ+vg5LpiUN/Pb8xf+zgo/qZfm70xnm1Nkp
wsO1YOKA/AWaXv8/FbWXdzNUJ6zNmJQ+FUv0TP+hV/+nTYndBgJqFle6vsg06g1bPRJt0fYtsg2D
resUqh7yg0bhtxUW+v/hjcq2nXHk6R3INVxxy0ZYRKE/07SU6hXqS6VPTbEAnDZNuVrMt7xPQdki
tRQfFmvpB1nxrDdohvo68gDRSWXryidX/KxhHFbhhcNyP8wlftwtQggGnQ9eX5wqxnYmD4FhhIyE
EYb4d4qd5rtKs9matT2ax1RTMgrO2NaMnYb9yros78HRY1U9AkLeQWB+iSxrr76bK61A/0JnpZfW
dmS09je1Ue/KlcchKonG+Vk+iiP7ejmQyQ57HxbrY370/LylgOMnHqb0XnkfI2Z2FkV48lZyecAV
jyPu7jQzRlVHVvzEM8h0ijzkwLyhID5dLyjBU9KDPsTcAEBAjzCW+YodhZVxjSxCxCEsUzLcIpAg
gdKKLUYDB7hN9uwAGA1Kl96JtzSH9cpwJ1chVUKqD7yfA2pv+GrImztepYX5ZfEFQxmsPNL3WMBX
aG0oI8vP+BHouMIUYy+8/dCyhETLEh5Khjn9KFxAGSnx4aze6tVc3TBloIKWkDeiBCtFVNwhQ7FG
LkS7S+WDo9H1RHrYvDOvV6LCruSB+CtltHMDWhp92fWn4qI0PXCwAa9SwZnNkMc1DD08TIRLowoD
RqrSkDiTIsT+9J7gJMa471kZRVd7s9jSKS8Pv/ctvAJTzct6uCF30QIJViGzKckWrdeUx00dug7u
x8p6wyzUo1jKiQUHfnrGJwZC9iHvNg056Db337J9TmrUIlC/2tKtcviJNZsqH7ZkXyJw8KbhPP9T
Cg4qDmkIoKqrgcbXPLgDQdmn0+9o3o8N543ijEyFeYE4jrJ+w5mk6tHiJ5lgZnYOJeJB6gZAoNvQ
gp5NNHLWDC49UBFfnj0EphPZhMP5Ipvr+26lheuyboUKBOlvVxuXbOAmRJY0q3mEFuV3pFCP8xKA
8qsgvxTJk4b2WlDKLpkCZsy8vmftnF6cVE3UEp9ozeOHcjMmACQuKgfSZ9j3RYsdsW1uPjKPE/k7
1BkPq/mQNtPWLN2f0YbHPPNo6YvC5/JSeoYIqp/BRJJj4oXAIWLvPuhsnCLKa2ZMWArNJgmT5gAe
wdFNWeFlEOnZApEUtIfrt868BhIA90XEWB5pugTByUKOpThZZMd0Hw2iVtlSI0GZYQR4zvqLLOWp
I+sHzvNAb+keZ2HbQCb4uNt4+Fhx1RrtiltXcT6YCPoqFP84g+cl05xe5BmzcCjevTB1v8FanrmF
917VN4bUqEdAveVXMkZsWM6lkq45JJKQZSveK0EpjDSShgPgcFKqzd3FVjYtlJbmTr0TKGB5wJC6
eLTX42oYlLzvNoU28eK78PiLwP16zL6p4Rqf/4WBxEsLvepGDv4phYzMM1NY/E4ti9///PBwTbVj
Mwl8OO6eSSU5CRKe3dhr375y8kKY63vw4R/zV00yIfSM0BV/NFZ7dOCJuU+Qkoo5QFnhEe7zBaKV
qmjWM2AMKeNj2Kxp1X0jtrjwmpzg/Z3MRJclIRcvKXwZ/OL82PVeNE7gC76zvqjtbJLmxLcofjvB
MbTZGfyDhJnC3APFnYQPhTPoT/nq9e3pGBFNIH7JhVSnYVdW38O/m2VzzWUVJae6uqhqm1hytE4k
t/lQGf8Mb1ZqMvBenQ88rtrXhFQqSZBIH7YPAl1UT2neuSmtO8EXT7a/TWtxvjQcEcim7707PSDD
Qp/TtlFwsGU1+zzQG6XO/+BTge6aa9aGK/6M7bCVQEizpWXFV9pHC0oLKuLf6HXMvqS/TlRwLtvI
sLJKPL7aSOGEhygsaYiQgZM0E48Ee0vqJhDEpRKXR++OucKkJRGJzN+4XfvzysAjaYwLVLttwkGM
A2GHyYCFT+g+coxBXvEMnXxXbBHgeY5WqtGX+lItPd5fkb9qSmC29Rxq/sCtO73wgtGhKYzFFL3B
gsCTu6XG2wGwkqmAlbtF7KQhBgboyfK5ljNcXR/f73GbMltjjGuCx9Ek3WY6QpJFx85HuKZvEjhE
OXKrYYBiZUG75B9xGQvaCZW9N24M/16jD8E67ngY6JU1GSYtYgrGv5B3TGuVbrxW4JEIDTk/8QTb
Tv3jGe05HZ1O4Z/qwOGATFHRBEAkGxk1RbKo9klZXPMAW5HNvmL+6DjdU8i6Mjawcw7jt8APhC86
XC1ufGpAq7b9bnWKbTDeihUeuINxO6xjoDxW9c2nzQQq40Bkpy+vseDHG3IPLnK0PX12qUOgRrOG
fG3WMg2UeTf5qxCOthZ18eMwv8H9nWvyXgGB4d0RGCyZPB9BOJZ4qHDy5BOpVLsB31vGjBEtohvU
NMR55Fpux4ohJInuHTp6wod34zMirVwG/2wHYPCzt3cpBvy2DlbV2qlOlM4bc7m/XR/fAeUNkn7r
NNuNmlpNSuFnmLeqRyssW8tgwS4L5SO4mD2tdZ+z9W02dgILUCMpEv0bpRB7LNVJjAkVGSITTHos
y0BcSWQBgezQrvp/GCDu1TdEvNR/9ib4Pib1q9nuiijFMBsEU/iMSnm81cR7jItSqKJz5jbC4N0H
UBX3ULFWrp3kwZQYmo5dlS7q6xa1WtS0sHVdn/9jxf1LngJG8rQgmB1SssirusbVPSOzc5aAkrWK
RPqf1tdiUGZ/1VsLodspIvLg6tYDDNmIo0gjOkh4oA4T9qdiLywYPvUdd4b5WIpjAOZBZccGl+Rz
/y4amcZAri4MM1I1u+UQtGlLf83fQG4vtxizZkOgxDAC9sGUdIkitjWvwS525KSWPMFK/AeOv8gj
K37lH4nuA8VumQKU2XFxMW3ALHz5Uyzczg0hDGuGRwpk1ZMLrhV5NuTJam0Vjb24a1ooh7JWkgB9
+vxbBm6oL13JfOsMQpcWjAbIjEt6adQ8/Oo9ZjdTMkns41ry4tOHbX9rGgU44q5HS5k4ClISu+D1
2/Y03KHb2m9/o/nx3ug3eG5QTdZ25fmfQUJOEpYnvDpARI8yotXlCrZhXRTPukbPfR9oyZdoYGmy
WyWNOI741qHSb8CeJE5HOH36Vm0OxsJPnQUD6lGrznED62DxIki3yo23dofAtISgeh/bvZ39K0ln
Yvv1yMdbedZIm6ZS3raxIfXRcgotXkzr+QtXeFqITW7JAKALv+0jD1jhMEf42Qy0EcJe1NLMQkDK
doh5t0xGfWXFAJEN4FJce/XdOXvVuogYzqpjW2frEfnyMs6iX8Y97YmfOtZ+dNxlA/XE4xRwCide
hjT8m9ARQtjcbGHsqCb59IaxH0OkTeD3lM5GJqE9VDpYNJIjzhLg85kd0x9VxMU6mSXduFTd0QWS
cyOzS9g7S1+wIq6b/vpHLmPhRYaUjoIO9dcuU3OnKoKUXem+Xu5LrzF6KLhcc4+JE9/z4yKeC6HC
gedR5qzTFmny67wQiluCLP7DzQVXVgqvxPXu51kxVKdVNr/JiJvZlaKl229oFNfxbT0haae+c2X6
BwJ/gCQchXKdq42LbB4JVxV1EY+ZEEiIlEUBftcbfdm4lKAtt7W9xnS8+oMF7xeiDqhUCYjEoKzk
16N9y6te+mnZX9/MXEotQksiT0VUW2O+c+T+Kj1MiDjxmmQuQjoHa4y8FZU1J4UYqA3JJd++bezz
jACoM4167owmnJfQeMiEXQtr0+ovxqkpL6Td7nr7nkt6WY1LjsECQ6+MS71lDzVFypzg6HqCTDfo
svxvDzeg8ej7EhCnxfboqLz8J+uPQH6l+/CP7vggmrP4hrWrBpwQ+sAssjVhsUxKlWJblDKxsf8r
VSrYW6XefliPoVEPslIPQbAQkAQ4i+iMCYqv58C3NyU3TO/Qbg+0XEq3g5kTfOr8+/6JhY4kERFw
jS6oUstf0J19oA/nENvCEid6jxTnU3EbjyWoYvh1WDcBZmFnx7K26Z5JNpbFntbbIo3i6y6Dr6Tv
RRAyg4u0Mf5pMaVRrFXVEjL093FTdIE3z/PLUH6arQ7aLK+UFi7RegqRMztZN+Kw+0bCjN2+Zh2s
DTfl3/Kq9N1HWudE/66SkDilwD0aXx8eKeErfMsW7Ozu2kNCZFHdsfor3dKR1pMdqjFtyTArmvcX
lTiIFOGWjsitQ+yCFggJhL1dLGOdQwPPydcOpE/7Z3iSnAIq6QyDdoi62ajANceRPdoqhf8IhxjJ
vM4nB92/aGRuoEiCjXLO9nTD46sJ/6VmEA3RJ2F0/dDrZ4tjCdd2B/pYL0Kmkaua9legpAqY70Cg
Px9++7pnoFzpL0zRI2u4G/CZ5eIqUDhCKkDzI3T4kz3we+ae7qofzPSwm/dAfnVdvM8G8998FkJK
GoYNcZv35vhySse/2ss2LNAc6yx4LFco5jpiRrrAI+vhFtkOrSw2Cy/DVPn3Ed7DQRo3h46C28e4
ab3TVHVZGysqPKsygsXVIMxXbypg/XetxzaPpuZxdwUavLcVnN+j95z1buVOdt60SSUC4V1Ht/vH
gJyiAZTXGj8FMjlsCQYX/vbqTaC9Y/ySFcc/yuQ2MNrgqrgrYKnxiTXsCF8s5kKrgbeoUzWtpIoo
66VZy6BLA4YSF9HhT5RoA4Dp09TDaTfHA8NXhOt53NA58uazaZ1qtW5A0aHJSoxGoOkiFhHyCAd1
E9fhqGqa7M/3xNU1Jd1cQz2QBCq0H8qEkeizEO5rggCBXKnVwJdGa/nUjRs3YPfC7ag39SwSEnHf
9cGV4fT8WlzT6uZCM8gVPKK8OD/UshbUp22rwFdhi+ZVInicdzyjM5ehhgW/uBsprzmLI6sn3p6Q
Ug2YnnqB0zoD7ykzjS77GFR7TVyhmKia6N85pvHzuBGg9SNOD1z2JjPm6lbYTdV5xbghR4/msipA
AmOdIFxh5ZQNJ5Kpz6Vywkiw20LbHERgJRdAaj1A+mAU26OskkFU8i8T33n5xKxZblefVxtceagQ
ubDOlW8SqU2XvUSsgoCrE26mcq3nWochmP3C3yQ8TbkMlpwjxXq9lMx99inIw7KOPrKyXrfKOF5l
Oenm/3cm3pyO205iJdp2A39ulEQq2vQ00Y5D3Clb2ftXlmpDiQK9x6LGmXw8K8PGkY3+QtDfEFY+
03QYn+lRyQRe6++As6cRir2rYwQ0vLEW1SAI23S6pbbtzML7BHc29b3t6TlqgRGTMXxe2MyQ0SBs
0I29uEy6VpuKtHO4Zh/QT4nIy0tjxY4K2WuDnjazaK6g6vMsJ3oHu4M0PhCKcVN81CVgBtXq1GSe
Zm+AmgF1vWMLqIL6imgnIuQrdt44JIFN4zoAQfsVNzO0Rl8S8wbY0tvagul85e5n6Ei+Jo5YGpo+
ftlUgAgAQlL3ChN+mhP+p+qIjKwHOJw6dlRI8KPPrVJgmH18dwwy55Zd81jt9fENn73HPAyrZy1z
HEQ1peq7/7XbQM198kt0IESBT+Qezx6yK6ggsTPM8O98P8m+BzlWezSU0x5y46Bj83/Z2grmoyz1
k1Zuh7nPlD97ERb8dBHUmgFHQ3LEPYU7CFHs6QDQFwK7TL1Y6EeUUYaX/ZPL5mDpodBVxxuTJAKn
t/PH1VoDTOZm1YVMsmOOY5QXlhe1h+DuTtIRbxPf19Si+1TKB0lbB7rmCG8aCjyTkXu9H6qauEiI
Od4owRPD3B98bSAxGpe3VoEkefz7m7Mi/E70V0Hh7KUeexl/4r6ktN6RWH32x88kO1WUUDOlmb75
KMVOYWnPCiO7jgyvU0u3hGlb3yOkAkbPPsWmF9gdW31OIJ0GetqcVY+M9XhM+X+9JTDARJuQ4S0k
y5kkqbarni0WpK+5pFYJhm/uuPTzBZsCIkTYnq9If4Axcg1Cv4NkIXBkFuBnBMYJqcwD+esA+0+0
4/+LEmZPMxZdOO4j5CGfmrE2jCk6kNpKCfztXneJ4+RzPFsY25iTXNUUYNO0tvmsJNyHcwrUNOW8
2PiTdG9dAtRnp82jGcl9W6vrBAKHCxAnHe5d2afgolOP9tBwUne4KKjDZkko1RNN3bwyN5urxflA
C3Nm4/aCJKa0lkXcS7NyE1ejUjZDcja4uuJRFXMKtKvLBgD5Nbialxnh8PBnIA2UHiOz+I+M14EO
A2rAPfIKBWp6qZHX0xJ/8Ody+vX8Nq4Trzo44c6G+TyS5q4sDQ9x4DkNa2T6RRV2mUDjVdc71l0O
XfnogplNdRKuSFQT59eaDGdOgO7xOUBQ8lWov/3IQU8OVIqQFOvCgi3cve4ef1zGWL1+JFr7LXaA
1APjt4PvulZDtlvlkfWr/t5Rlraky31pwLFrY52AH2qkyCbrFNDdk7yK/sX9M+Ildh4TOufpZpV9
R7VxV4WUoV0uQmVCWpn1jKDrmAa4ej6EXAWHwJv8XRKH0zCtH2RrroVrtC89yeCyYg8FrDcVDmMo
aCK3luqZtSvWDz1Zx5NGVpP31LtwjuHRCrDxdSdP8y3tuw6JJUohUGOT8DaPfA807ZcRRUSP5feA
mS3vdYIdbZo9aHo7NUhUYcDyK9LLhb2rQfRur4AdvTrbKORT3IJJcSmp4LCJ7KCP720t3oSNerJA
EP2GnvyiqUFDDuJhBS8WhjGnZd8r6XCj3H/0CSaPYT4wR+1l/2a5R/gI1bvvcA+l/RkplZeG0tA7
4p6CfLc/Vg836O+S2q8OXKHKnnG2jl/V2JpWB+AMb0XMIvaCDBF7pGooN7Wq3Ht3aeTJWCsUUUcT
YAi6J0TzJI1nMmoM/1CDscbl1O2omF7uoLr6+BQ1iqtixy23EdJNSYE8BpV77rOumZjoT0VVkoFI
ASbKwdiC11b5PDDPeL02FcVA8fhLQLMe+SDiYvK0f4Ec85TyWm23bfDnFhiRxgF5DeTlJhbMP2w0
aEyHZj1vO9VXVtQQOi3YluTvqvnjZJgFhETo4scABeiMfgHPW1WezMchLbkTbM+eb+FVhSoyBl+g
ByeKna/yzNn9gpNS1BGU6sfcuqaKpi43unW8/kz/6tLXyoYjSFHu5d6vefoWm+220+bTGkbyQm1R
GWWBspuw3i5Lo1kCHEj+qFbFLgeVNKKKBHOg98rsuiwb0WcI1YOAPCPao4ZDUjJTG0n7jFUD2SRi
kUt3Pjb8hYYQ6x22KiouuT5MDzP1zweLgMHww50Hr0xH3pjHamov+23m0kr5BrM1IFEHNHs2aS87
55Jrmz/ftwBkG+NdhbF58hXAmqyJG0iHEOei77YKXUa2XvE6JDSfIgTzNs+3kLI4uVWaB8IsFA/F
FYKmRn6J8zCIaaKY6yo2Uwj0WeI8fQJfviymdWxpK1RqA++Rdo+jVkjgquqMSb7QkUaWiSy7EJcE
HC7gKF5Hadhnp+dZ81XMzTLfqLM2aNKLk/8lYmFWJ9EL5IOxXsebq9N1+ScstSe20N955G5c4iZW
/ndjWD1reKYwXmhbfuIbiQqpNOmZY7OurfUqij8wQA1+yRib3l1cruHXQcn6oRpKJW1ZZtA4KMUd
pTu3EFe1F2XatCpNgb/af+JlFdqbYu5LpNa+DgPpfdFTpHM5HMRaTTO09ThPKCPBAMyeNgooQMoq
DlKH1jE+gHDOqpc9GnPCGESiayPzutc1rNx6RrnPlHmcrY0uaxQV3OUtLifLcrj5L8S+gKmpRfMz
Mw21KfjOe63H2Rv0HFvXWexE0zdbxazBXJHgaRhpTzEaqNDB2OT4RMRQkZIY+oak2rxRnebUanzV
BGp/4DPnGBDMrcdLPKytMo5qTEJJNaGS6b57xByjg3HXyEUvwLbhNmrJu7eAfm9nvqizdpGCAmFz
GjmuJX/Pv8PKakc7a9bERSufB16HK3WlQc4Y6cVeosvS1nOy4H+9ZKj9Tr6rTtmoTuA32KrIaZ4a
+dSdvXfl5UqXm46K9MsbKqM2Hs0w6NmhH+15XdJh6RWh1f4uHldKIWmIHtbL/SJop9Lnb8TxnVMv
QGe/EnLOTLUeiHd8pCqjkxsRf4Y2p9/fOFxHzcRaArgtiyEUkddkQ4BLK28C/vuggQ1gV8PuOiyG
44Hp3xwFeXI7422xhP5SLjzY3njdE5q7pK1hLUaK8NB1d1h3F/GNlIls9OnbIAHdyddZRvP2yT2e
+W3ZCv29GuchjA5RelyTL36kzS5SW+r1w8A7JPVfZw/PKKY7POT3GjtNdMXosAUG9N0ZmKoin16P
j9BtS3zs9vsXx83l9PMddq/2W53pgSsEBEio5IaNat/KkfZ0PaN6vgBnBdzXwjXD0xQHdjCkoQD5
WycWLPTxyoLnWtBSoweFBEc81moNPoAxV0pmbZHmWOuv6ekmRJ2I1EsFgpV+GFQ7FLu5FhuqB90d
AxjhP46ShLeL56ZVA9EgpNVrSvmUtn+Wz3S2Y02Bg6GfOc0H7U25BH1tI5Ii02TvdoWoMsM6F3gw
dDmWpQmA52S3FdZNKAQAwbYfXZUF+cUGCMNeiJSOyACc4fODPD7AS3y3NpaFC6rUz03tTuRUVHMb
KAptpMNfHz+UfInP7YWk09UEprcioIPFe8AkAIriNMCebHjaBpz/Dh4R4lIR5TecAlH9bCM2D2oX
jEIzD+3E1bxTsM5Y7DUDD9LKJjO8QC7h8EvnSFu+fJmFbb5bJagWh8iBHhCR0c4Kb+mirapt8NMZ
Rdt1kd6Qrz6Mzp2YSO3tgOpgul6MMdY5MIIkFT9eS9yVA3ib7a+u7Q6khoU3aJol8vo7DSmlcIXH
603Z86B6kyjLPh94L7czK0XYH5LLl998Gpwc8s/QfpZwDAnuWGNAvNCUUhDPZACQsSs9S7aJ2sbG
lDLVJBKeyq/nrsei8weVWO44YICG1hKehy6AMApK2PGYIzWrX76mVHrs6bLao/iEjqE6tJ/soxgd
ZzCHxgkxffkkj/E33JBV7I5z4JWiuBNGH0FDsTuIbyRBioCW2BWTmZ8/4PE2H7M8BOsvoWkCKR5p
vdtURIXZrclgNiEQJGeO2ypB9DQ5mtT+yqPFeP51e4tlTePf13EEpxnPZV1SQ0fCg7mUwC3uuonl
b+GRhUDdWaaPX1xd6q8IK1jm+I8m7KNsesHeJhUaWsrdGtaQQRfTjccCMVXFLkUUhOQuItFGzL0K
R8oKIe3IKPGK4Ywyc3xv4CYrGzUQfcS8578Wz0IozaK6AQ5bnKnbqbTF5lJNGp0b1tuQ3zp9PuNN
wdlSLZ8q/S1SI7yWrbVkVTYpOWJEYdJ+LNb+sRlyUUfkdbG12FGTL5WSMrTvwiYE7nw3GO2TwhNj
7cJfGJzudXmjlhD0VzHriCSMBUQGQgH/zyYdgpZgLRFmAVnT7C72HjfPVuaelzvbtvCYaXRVJx1I
jtYC8J3eb+GXW4ddSNqbMO20u9yzMv89MnagPHJnZR9QuyrYj9U9Wd47DgDvFWJDe9A4OZS4kyeO
3HvUpmn9hkC6QM+wK4N1C6jw+zQ13GOCeYjoM7ECyjMPP8jLl31oUHW+29Uzm7VCQrK2u7/JWp7Z
SvxJ9n7Qd5j3uqlD6eguvNzuddIVXoGEusvR8UaWmirVgAaSRU0m4MAeZ7HqdR0cUIlF6UUkXAAQ
ay1Z7mbP7Kb+AM5EurJtCIO1vM2GjC5xCVPmQTnbELpRcHXxJoQdKG2TiB0ujTYn+3tzTOYZccaG
b51Be1FsmqNzzBxJunNnT1MI52vtdxoTfOQQRA7fhyDU8bEpmkMt6XDijGxx3edW5V4Xfp3d8uEC
kd5DRAz/zkmA7WAyRd2LIeo+0mIyqjP4JE0joTao4d4965fMThLOwWU6TOTxSsaNon6KwtS4OAez
yMVECL2Vqiue1aUvSiZremxYfO4X9ztzV93hY58rmdhd8JaTurmH/iUn+BBxsstJNH74dLqHEGl2
2gG+P3r/XCh9YC+N8WS5ehvE4eJ8RlNYXwmWiTIcd/XOF2OwIWn2tzaOYCmmBMUS5DNo1G0RUWQv
Axd5L5tL3BzznolqreR2pjsI1N885brJeOShc2TLgYmOu+KTVRhUZyf+IpSNZXJiL7TVlsQRj9B2
AntImXtvlsdBhcVgSm5PHqZZGMUb5HLeKLDhNnr9ZKA7a0UcWTJeltMsC+EBaxVVuhHmGyp+zS2J
fLz4rJ959VqgCLi7ZiNVM/H+iOIm19d8Q8UN06/FAnCQQdnmxiNlTqJ9MHz1tpP4apOZOcbuubyr
Gg4odPTut065Eiu5TuhcxtOSSOqfani0U1ck3s/CDb18VzsT49DbP78LW+ElFfWUx8gz753T7nxp
CC5C5yRRZcDjhE+7L5PXclXHAggq/fHRRYGS46wMJkt2Rw06wtuTaZCDSNeBOX66nobsQ+yieUVd
gWG8ZQZynpb4Vox53xxFGkxHDwDaGQhKJxMUhb1iDi44dDKJX64ETatEDG79/RNGzAuSQugyXEHP
mfGO8kSBbIhSdyPvljKkGIk/x6SxwpmeWDh2pMze5umhqzuHTB/ZQisOI3YgyAnOb3Q8YDDRQSiu
faqe49ewecXY6ekFNpYe20NXgKN4VDrPJEKP1OtBH5P2FqQ2vwG9uEp/7A2sqTKvVG8O9kJNeOHM
XW3RMGRQaufKB5e8KvK3uBO0DjAmH5RBhOJivI5F0DHnLQc6FL+y5oYeacofdp6d1ZeLzbljeisf
dy6ma/GrE0tTquDTWE2bZjmDEsL5SEa0aqW+nSduy0ZcncH76bVebdfThjTcxYnrYXQAn/vSovAK
zIP8ERTA+eCDp9LUyoWf9uv6iqJwVu1EgjVceKBk3HQXrOid7BE6tD7nN5uSGFUogYFynDJGefYR
3ZC+EKGtX5RiJ5oh03SzGgoKOFH/L+lMWd88SIozNioqTeYBp8Di222YlWZJT6XfkVHiipfE5fiB
CLNXbaMynC+oYWtgbVDaPMiNdJ8QYt0U0IT6lA+6sEGLrTrc31d6Ec7jrf2pwMnaAjpe731o5hgg
tkjHtL3x08QfAZRgccEw0Cn7IKIoro/DakaYXbrDatuNezgltf8D/04TgNhcyRetJtudO5tY/IRQ
Xcm7lcRoe7++LyssCtVXE+bn0aTtSJEnO4tJwBgeSlsKH0WzpDUjBH37yT81Rqrdm3x07JZD6DS+
cHIJqervhhozbFACMsIXfVpiIktCZlzO1FgC2MRA+C9CLNh0Hi4ZokBmViLFKgpkW/JXvqC1x8+G
uaoZKN2b2j3dAOVwnHcjbjgta8SPVaxDMCq9JqYCr7ccCmlhTuHkxV3YeDLduZZdXJYP6ADajICc
3Tk+CeZKMAbJZYRt3FfLeYASGGmu4tzeAkdflu454a0+kZEDHdKvRMnpv6sBJ33ZkjbrdJmHhPAp
Eb9/xlRlbANwpwN9fGT4jBxuEOoMJAHNHy1Je/UWaUOmnFhf7l34XGNKPxb6ABguvIm39p4A2IMM
9JttHZVY6n9eTYcRw5A08Pik54BbLEr97jeT8bPw+Q6ZRjiJL/kgiuK37oRjaVVDKWBKlh/B50wN
DCBPYhOw7dMg38DRIm5glH01bizykRkum1WrQBAjVYHascAqZmZYJ0RNic6HzHjPp3GB6jbt5ePc
ZLg/kaB2ltLudIJWzmrN0HYfdl9O8/L72JyiBz3fGw3UObBsRzd9X8gUavQEq9yhzCiLi5wninCV
8HxBdFyuxwP6l+9AP9M0S5AVbjbTCbppemWdJwj4coG8DIMQ4sq8ceJVUUS6hLllWlWCvYflM+6B
RhNjRWMwG9ZzFPW51o0X7D0m5AYYgQvo8TlIMpdwglhT9b1Ppb//ejwrauNLIfwFkLu90GHDNcyD
CEFvMO77fdLQhUcXAOt/dCDU6R5fIyOGWtVLwP1z8CaNY5R92yYu9TnFC1s7Xu8imGjnXI7yIm4H
/A4lqtzy7W8BImg3wb4f6Zc58/+eRgX5hSUl0IGqJ+Zzy96V24En8sfTztK+hWEtn6+/x17LqBVC
n4odL6QduAMCIcSgt+ODZJMYXgVAYfQWZSMdhQ1RZao+b1Vlh9lu0Z0OK3FyqaFXl9TpueJ7UQ5b
SGtX/+uQWAgGaz3/OdzHteamK/mP/VT83m7vQs44JWu+hv/X9gHO4qUX9rlGug+Nd/ewd5ot0hm2
u5NDepxINBebzNYxZFKHWI6qz0+KA6ZPpikBRJxBD12xcTDZtZCp0PyVFDAfTPyuiPz9K/G4TGSx
5njdvZDZOofuBbyxo/LvTNPXlEenRpB9E2knzLdAIR+w9Un3IJ8PFjaiUlxpK1QBsHCyk32Yuazv
tAryTMvTrp/hTG88gp14Qfara24RJSrjx+/Pludtmzvr4bYrWKiRymf33Ti3VOrlyac/pBUKPbtC
u0Oj9oXiQEkb4WZw8PCiFDhvJU+7VymZS0HmC8Smd26DLTgj0zligOGJi/3TnKwt/PnROGDY1Tpw
Fh9x23Ft7RxA/AOmit2is3OFFNqQHn8E3F/w7ioNBJ/xYZWiQouiftLAh2LWxRLdnio7gh26357W
gsDxoPreDnIoXi7Bj1/N8HOg5sfUQJXnyBw4qXTqLxb8+k7uV6juMQxB/q/eXl4EI5ul0WOSbvFy
DbENzUNUquaW+FFRVRuCoUloZomWeWenibdDrZ5sDW9dNi4HtFX/h3GToP2+jMkrduc4PRo8wMrA
2h4dOumAowBJ9UF/z9bvGdQFICmgw/R+e4in98yTNgKQVLa4B2XxX/4rP0MeI4nN86VPET8VTZSW
JT8V8IGY6uKEO6c9VEnchVtMsTqJFQqmdQDs+MdAUr9stX1WZydBeSP0TzF+rDPlgXooI9xyiDts
m6rrSyJ7Cgr5UnBbKKOF0Ut+jG/o/BoGrMuQ/LlM2gfWsocme9chWWM9avuB/s2IiF345TgNCJyy
jDkPRfbQ4fclDIPE7ZTmrT0N/Cte8RXC897xf4WL/fgZ4PLezn1ex/+bEsuU7ulJkcGWMpnwO3XX
fngnD78JSdAfVBcjcdyT8eUwF5juaA3EJiRNMTnDDbCVk9y8Jnzufix2ScUqBz0/BcMyWCeeL9j6
gy7+4WHCWtBP0rMyxbxhigM44Qop/GIFbNXhxK3W/JoEhtLWG7H+RKHlkEXzjVVivGNUuWzCFjLd
qOCzqcMbC8gAfT/d4EdHpyiZyOkuHk3Ejjx7uSkq0GenVQSP6mbafBCaiGbn97nlwXnKrY7oKizR
knRQjGPJUjgaGyHezd+YK2gUqAuGdEQcLVHYkLGfbV5i0SJO+bODNlgGmLq1uCbWoX+oXJ856Iss
nV3M42h0RZD8wGjrziHsi+Y50SeB9GlMgU9avuOqBsotp/XLZ4qkmkIdLqUGv6BsvzOb4y9BCEr1
x8qZFdYsmdXluYra28yoYqVnqwj0KH7NugjiBjq6e9vJeepPtqMdkW29vLH7inwpDl7B2eN93wIv
tswXE7BHbSQMgnOyXPNNsfQnkxvYRVJhaSiKe7UjGd6Kx7lLjSkUCYyxaxXfN+swGOP8Vxn1P93H
DGeUx3g/DoYMhzslQc8sYat0sbzKQH0BdGctBvp1wHrSW+TM3tAGEdnCqG35KHAIft93TMzkdtvS
iHBjP05DO9UMHIWhEiX4HFgsTdJgQ1gKIJvAw3UDXv7CSeFIEcQXOsOaG0A4+Z2b4pkzdznw0II0
eGy1T2UPQD56dshKo3zQCKAPSvip4O3QBLLvSFBhr4M4B2rqFx553eLQ+tdE7kPBgPLnlYbUUcXp
vppa8QWw1I2bg1VLrdnczLMPrON0Kroh4yvAXJ+EpKo5kTgLw+hm0MGjGos454x5+hZ1BYrFfAUq
Lz+4Er40kCAY8CJxRlSAD5939R0Uzycs54pP3TwrmEmd6luXpavDPO8P7wWulpewv7rIwvyTRR9X
Z+g3nKCJaPYgsfkSWYFBYGUn5IYdMCKaQegavQc74k8KL9O2gnxwMJcaxtf0xY5vmBSl3ElGuClC
yWdXrQFcl4Fr/nclHsFL6IenZWx7RU8Z9WYED5sNuOFxK3QBT5cS+WuQmJ/i1ve0tsRlcjEew2b2
b/TJ31TsEsq9ThIqp0mYKo38gvbvjgFr8clZ7P80dhkUgV/0VPsw/9TBg31q2iqJ13BuOkrz5g84
wP9k7umdNK9hFrIZ1A53xNJDxpllyGKI8o+vQ6eDlsSoGNA7awgRubfbSftUXJEdp/bpxLI/C4bR
JqP3+kGXdZ/WO/Jcg1TzbF7KjDLF0/290uwSURCTyOsZ2WK+L/cnYiomK4nH8pEr3/w/bIHfohpX
zcJnPRVDM7bt7lI9BKi5rNUegHsVgqJhnFOG9bq68Bmjpq7A//qdrqD1/CGdzR+lwEfJ+k+D+a1B
1SFu8JPvmHpVUtNVfu/NztdTwd20tcrZc92ujz4VhMnTUnOjOge9QGv49OBY08HkKy/TcDdtlvWF
7EO5BNHvm+sRpTZploycsaXpLSp/1J4s5wuLNCZYI+Qp+1NpSWjD2jjXwWDd32XaCCwM1WEsOW1m
gprBmcJIu4oVZzlCyFCPxvywUapChH5IaXuFcMdgtMVctnKCHM0Wp8F4rWrAHJcTUs2YSymdGIwi
YEHWhQIvCy7VKWrFt/nSlhWhfHeCnO8rLro0nmhA1ESEH9a7EaZwypjylEDa6b8nqM5PHH3WBNYu
N20zwEUUVVsypElpsJs6XJBPJDlOlWp7hc/Bw/QMNdJ+0knueBmRp2XVxjxwHZy1MvU4fflbWdO/
zel6WBPKQFIsc49SikCU6FFU5whPBGpZ6GCckcQTUmwNncsioxvB8Pjgl2R7N3gbgg1LyDVj6TEg
Oc3wxTzmP0MkqsS0Kmec0XlE3kjJBDRzpxmqgdBOgJpoEoBIaoW37y47qgfylMLJLJpCBMxoByEy
G+QEp3baTc3tmgoT9FMEAh8tKgg6EyrQj3AbdQxLhD2rh8G62XFkAl5O2YWBo3kb7ZEe7aefDDJt
roQpCdGRGybT2oZeK9hEHHuWe/VJhj8c+2WGYQ4bm+6YsRJCKUOuHUmzH/aMtP2Bhsr5wl9oZsuf
ykOtbNhFmAyHqawxRzwbF/IGZLBOiKc4sI3LufuJ4xVJhVO9LOiAkdHO2AT1aHEYcUFPQH3X2lPA
Nh7rz65boaKWL6O1vwhmGys+cqTUHZ0TJq2HvR34HUrxduAU4LlhUih47dVfmSksC8vMMfQQmT0Z
4VxS/CVdLclHaOIHdzU19qLTHuEkFMzAVPst9gZXL5rIUZUi8Lj8ibG5BRfzwkaQg8M8zh0F+Giw
lC7l7brNJli7kTHcTnst/AqYRSUR4andKb8dN++69PLSmBkdKo8Enxe6RNfqb1ceeqHtcj4GOS8i
Ez+YxME/EBZDecro38sO7XSH+pdAzaOGPMt9K5rO6Wu9bvxdhLEOyOyuB8cAtHcxgjHoxQo3Il9w
7sa400Az5ZFU4AvkyHB3iNOIANTQ09oZBG83zwiHMuqH2W66bqE2JE85ZIYVcVpKReBosUO3Rmsx
nutUOLUCkrjWVsT9MnyYaqagmQS+NbqGYoBqFGQkxsAq0cfg3PURndxmFlMwtqcsKQboocje+hAs
2I9Jqrtk9ABAvtYxY0vRGHktava/8QOhSBz099YFANtP20ADNc4vUXPL4ci8AaVXGhueooIcXPoY
IW4rjjJQbfwTPEcniheqfLFSLNoTiQDKNs6vDxz/UhO4GvAIsxIROlSPdIiRm2INt3T9VBQ5tjP1
Js7nhZIBOCSRLFpBP1Sgxve2WZ4G1v3l7p3h90oOFNZSl1tAATd+892Bm/OTdgc6O30/VT4+Dl7F
5kKDJkiX8DJ4GU9aaaHNyDAFEmZ/LdSvlXaKvhyHAJ0jzYkMFpx6aNAzR2A7p1c8ABrNL81ZABI+
m7T1rpVZgPMX2/GtXxvk8zdmGSkEobk7wECpo5k4pdygE8wFeyp07GNBgisjQB7agnoHlYn3vpgE
3Ar2pEhf2Doe6G7jbjt9o0muDdw7lm6gZYVOTSXNKl550tNnOjHgDaI7IR8JEH9AwX9AIc4bnG+M
PqFidB+bFcGHpSQjD94fOXDhwjnuJnAqfPASqCzuJyWQbKCiccYdZEQOXKxaDcxEZyccFAdRvOBB
tbUB1mX23QJAuFXi79LB26/Q3HP+JpyUuhFArzYoqMgm6Dh6fifpbEQvVpcJE6Epk77hz7fwr7OV
n4oX4FqY7hqCgjR0bQNLBM9Po8xakhe7Z/whHMSKzcKLf6B+j+kycb/A9+ODgrsvZEJSXDk5wcnC
PWvb5dC4BDZFl7ROD2BuUnBdPjfX5Q8QF7yFSFfQ200Sz2CG3TaItXDS3941+AVXstzLRbAvNdMm
EFqZ4u53UQMjrgeQ1McAvD6orTb9ucM1ZhbvidgGP2p8/kI3sYNr0Z3V4ZoI+DYdWn9rIcCY0qRI
r9i2fPhKbCe+ZPl57u3b18fM8D46diwGJSzlPvEDXIGF/oQwXApzlZ/+ykqixLNmtvxi+t7pHJW1
PjqmDmy3OKDrCvyLkvA2Ypq0t12wNEthjAP0HOwvwSvxPEBCYqe8NwC7rmiKh/5DJdQba37zB3va
60gsuC3kH3lhDUU7qquXHri6zyoOSWon8rDuVPGd2UF1KPMYcbdTYWgPrplbqvH1Zi74h6H81QNb
ysxgkzCtLwThqOhLaRgijU/xBuoYbdrw5fpHx146k0OM6GGYcDiM36RUR8Qc5h6SpsygevQ4mqnT
04hunVrUxTrnkNx85cdZLxu0ekElCOF6MGdtGmtsthtjVPn6Lz0P/nAOMr2VFlypx5AXfsF1exDE
jnOYdIvDbGXSCePllTsNgx7Mn1iOgvWGjCZqqTrNb7PR+8gumgb9DELTfqzYhm0m/wGjzZzVnYLH
TCnXBwM//VZfalmlQKjrjAHtnFYkCPS2qCW7VzstcEAVh3/rMZeckvmBh+0rvt9P6j4aH4BZfW14
j6rHXp8hItMzWgXNRZb85goaMxRpArBFXh+18s4tO8rU0CVRSGZZSL7X376IVSIZMMohJE5zUe+s
iRtK/xfZTNPI18WL/3jChR5U8wOBAhYpCsxQixmOJKHKzNG1KKV1AIHjepGZxYHaogGugaVu8AIK
Rbj2TO8838CHx/9c8AudDtrA+Ooq53AXFZ68j9k5rUSv2vokHK+/O4FwXhQD+bNMVtCTrk+Nr/ji
DlM21Y9a2EBQx+sVdTqRdQ2DnR813H+72+d62H3GktVwgY66g7UgcBnEaaSwaYd9cLgF0Oa2sMSF
a2zqgmxWWucytB+rEGvfP9R2mZp9D+/j6WvAipISNxSZUhf6gV6wCkxu1C/DHgUDhhvGajOHNvLL
TPV9AeGLfHcxwH4rkWAJG7uCajOmXNp6xO+8QQvkk4W1iTYTYQaEhRPizVsvVivaWrintz6oa+us
MbkICCNXyg6dpzdHk1ZIazI7HRhusTyLcb/4LAR5UXZ9BY6zRArMobw0I7NIwtoD7VjwWq3iAYo2
cTh/jBPytzVFKNQI19/jTTV2bTR+exJbeJS0ja0uNWz8hwhxMsZlsfMQYU3Ahf0gshbJZqWfiLVH
jEHpFq7IYTfdwWkPRD2WlfPJyW164OB03ewwAUSZqwZC9oFCeRqfsV6UGiAPgyHaDkGTGu+k6xN7
KdVZGedIaXVnImn3j7FYptBUeD+8bG/4jxtNmtUSV8aGNTbh3XVAo8QiCXUVf/SMyZx73bCuvxAN
ddgEwns+2/2FvRevV/KUVIS0F5roOvbIh4PuBz93dJBbfZY1bOygEpsuqK78R/lrz2W5rL0PjNAI
wrqnqEdwcfw2Z/C8QeQt7IzIkONnR8bknMIhymNulhU6wy4wi78VxSv3H202NfQaYaq00iBcrXhk
F3kjBBm6ZdKyHMlGnCXaOwaT6n1RRrFnkSrWurCse6joZPEAgfyTxSs8N7dnQZRHSJ3H309CQQzm
tfrBj7gMtgcWcOxgLt3jjsx51VsjDwS1XTD65y6gka78nUGFqExvstYyhvi42ogIGQ0Mft+enKDm
0pN6LAa0u8KF/tf1+B9+bgQs06poIdKw7OVORbUVangchCp53QPWyXPL0dsbd/7uZy/UsmFCtwRg
9DpO6z+njFr5tFymTawv0nXSuY9ttnTgNkzoiY2X7NUkXO771sc57NdpSn3DAi+60GZ81v0qKiRf
yRsc/KUiTX6q44w3t5efodK9pL6eYbMg9kSjjau9BesOvh+MOUvnoQeebslQW9HMjUyvvnJuLc9f
4MN0izvmlKmHpGjZr/vBW+6aIVRmDc7hXsNpFS1qGLjSAH1fPPNTS11ljExc50+sMLx8WhXU7gDe
MWCy9V/QdKnGHGFqCyDtzruSz//C5VOKDGWbbaLGDkZDOpSlPlR8/ZpYp1mKkqGp3k9FP8OvbR8O
VD4N3t6DqO6BNQ6rbHA1zVSVXinYYLRzA/3HaVopFcA9dB3W0CzcQ049oBoLtx1kPuIrAliOfc7H
rsxLDfU/OP3toLg5QrJh+8JOwShO306kj03KECrSFGm4y4hu8iyUI7TExbAsEqqskgS1fbX+0HGW
Ga6tjMN4q+rtYfUlhwHUaTP32rwKzm/LepNTOlpo7vPoa8V3Pim5DHTVoaUZeH2vZpDYfsy6E0Pu
YxrQdi1qQD76btaZHDZP53IAc5G58FfPko1vPRnfCXvq0TMy0Op5NMNiPxop5BrJrDklU+JesyXt
PktaZdA0pRH7bwfzYYxpW4q5wkbQg8hQQW13IY9TZ1qrILZGyAk4KgteXxXyy7UasHonq4BGs92l
PLFg15/+eKbb1LXgHp1DvQ3XTS2jD3iWSJ5+JKZSaSazgNzc9L2iN6HDZ7gd5O6bcZRruLUS1wLy
TilRfD0HjXjRrPu0jCH4/aXoFvaR+WJbzCS+8NFLsgv3+tR5PES5r/SMmsAPVDmeIfr7LdQbwtwF
r2JDLhnOAiTGk/6XAjzyPkrYveJKQYW7ldD66/VfSO54rmlAvcoqhu6ALoifj2r5crj1rpXHNDe5
bl7CiG/Is8m6VcKPhiOt1CwTs4L7fLLnQOKa3hJP8TLZ0RXPURvCWegfJtA/g7rTWEOFcHKaSE2D
Ct+fKKkCKpXtWw2oeJqZ/I/pglGKqTgJ06D0CiaqC7gGWY83pGrYm1UKLKLyFnhzgN7cK6GhO1BD
nfnQb+5km6c4sS5thOaVcHrae4JSMnhJfbqBXyZg4LMnzrj26zkcIAHn1rC8yJ+z0tPeY6GgLMpA
T8YDoP1VDPUrQ+5MAmtdCfI5TK4syj4bFkaamAjSQsZrmWZAvBodkgUWVFPInEi1F5CNFesAgHJO
uuu0aa+x1xbZaIDfL8WQqFY0lnODh7ZXKMjpZBttVy58YJ8CiGmA3nQOKRlG2jBXk1QIvVdUUmD0
kZ0qeqJvYi0akQRRyjOKx4FbifJChwSfTlUjnjEROg1DsUwGNvSmKMPe+KrEzU7ErY7GQPSgV2DZ
NYud+vl2oLU6t7rVCX9JwYBeiY+4R6ntKMQnieEc4n6yzVX1OHrsxWPtxQ/Vm24Gsi6LZMyrxTgm
HmU1bS8Cii1ojmWB0G4QISo74Sk4pnWDcw0Vokcz7rYyLWkgrKi+rlcNjV3VX5LDnjtfxn1+nzs8
eV73MH7KAO8a+u/OESSPhohtnfda8jSBVLxiyfZyl8wRzNS29YAc5f+6tw3v/8h+Tlr1m7Lkm8/P
yPc2zL9mkpI0vZt2inSJDmXZUF6/PXqDpHdMJe2Fewu6NJ5peEiocXbhkyYBXjwi4KE0wLNDKXiR
ARDmwqyJwxpDphJQ+GkTGOI6+zKGlRECn6xx/KAzL3GXZavbAgerQ5mAF2tZG0URBB+uQ7kPWE0R
nUPEgg87ilWTcJ1tB+wpu/H0I/bm3BqFXkYke6R0A4v4YfvHzJGE4hBM1DpnVNEbGp/Iw0DLs8Ot
NbFXqyz0KTlOOJZKi9ayNrYtkr+UJYgAADTEQ116wFCDAFhR+O9Jmz3rHfWo5+j6jBdXPTKPc82b
kyqWkoENXhdHd+c72zp8VNDR26rXYwUf3TZ91kb7wNQOp6wMWuaizX8KQ3qcP4vWr78tSgmn8osy
PtN4zNb+kXSJ94Nw47GyW7nHreUhcZCnXGUof8Z4DCilfG4tUA6xs5TS+mJQTBmZly0VbmPXsZOk
AiSxxAn6ayPCfNahRBdA4x4TzyxqHhLqOPFifBPFrPWzumtj2odfm5k4pPbtrGNEfb58skMcp1u+
lIDLCnEKjdZ8pyaW0r0UJ7ngNp6BciwlUto5dS0L7G1S2pr8ahqXXIjt4Iy+ZRkyMC6wjNW3cwWG
IPyrkT+8SLenDojbUK+llygizeirzEnIdxlHt6DHtEVO0vnz1HO9aEt6dDg44NS1n8nJTIgOk0Az
5wO/nrliuM5/XTPWKkbr9I/1pnl5lxxdJY5yB7nodfQUHghPuhRzANK/fIVBFKQFykr+4wzbtS09
q7txASvFf38jfX0DdhLolHHE07B0M+cI+F6Q1dUUnwPKq8NiDMI/58bO2gGhx0Z1auLTEbkOTOyf
fvU2Cc98BfccfC16o8gHtgQ6laCc5iBOWWf4KU1WFR1lFs74JFG8jpVojoRsa1wgpy3PHZ7iY3Wu
tj+CbmZH0xEnuz929rDLiNPrOYvee6+dr1Dk0bhUTbKUemh5d6XLoBdLKYCXLiLhBDXdeJPp8Ceb
f4iP+noPjyB6LeIfenatgizQae1webpvSiHEPi0vh2O4+FnJjAjiQPShpHK79cqHCuwpY6lpwESE
bylkw4sOJ0D3H6o5gIffVxjyY6aa6uRkdLUn/geyy9P8wHeSnXcAzs/Bq+chZSuGyxcF7HYMOthc
W6a4lb4vek6/AKwbCn+yuk++MBu6aVyMmibZ434XxNpkzmlNA2o7VfG4uts6xNTXmyxI0nbeJ7ZV
7McIr/7+bl5Z7L5iJbxFuOX04RzoP1X44bg+ohliVQF2YX6bO7//S8r4IoLxMBzE73erYrO7pUj5
7qrJv/UpmexYaYzL01NaFTsQq4JOkBMWZ/1jWRZzv9f28x59vY24Rkm3yiJA44MDUPsNxkHN523o
D/HVccKdRp5lN9r0TorPNm2ho7IAMjDuxUgPa6EB+lIYNlJUnzO+JDofZeAAMQYgcGGvVWlRZLO3
heUpm/DpUdI60z18/f6wyZLIrrBCrqPM+hHDKXAW36FE1c7n2vDNo77m7II+G41bgEgyGimhPa6m
M/dMSctIQTYv+G1jp7Wyo/XZii/fl77L64ywNX63u8AalhCRhVJlIon6Q13UYYEwW7u91J/yeIU8
9PjbqrS8LpSlWutEh/M8N3VdT7B5eUf5jOTK5hIMX6WIEbYoiYCO5Ixhgka2C2HZKbEK0hqV3pZU
eEbTx8pVSVxaWiUlO7OW/S1SzRhy7S8Ab3hEN3+/XJfOdFPDOqDUtUM5ibrzCF/npHzQxB+ATnQ2
4JN4NQCaRGrpFwvYFDojm5RKUau2D4e97pl1oi+KG4flaIdZx8OazBVyPZD7PyvdYDp7qEasHm8S
/5PHdb9yX4JXPcej1uLCYHKSkGZ1xiLAXQ3qvRJL2I4cc8YDKIYVtLoexPBEx+vy7x0xFus+XhdR
fS11QgjW3uEfdh6LD9uv7tmqCGWh2WnFG+OTZgCCP25kVaPECKifh5bjL3K9hJP+alQ06eQfGc2x
DdUL/Cu/QiUc+j3lNsaHCeF0iPCVxbcG6Fllij7CvOItuCcR2PYgXkVeEqnr+7kujYHAHU+YFDkW
rRc50+xwn2UhNaIPkI5zeNzundrDGofG+vzFariPuFg2LQlhB7eqo8Ut3jy+pCwNMjNI20EdIyle
an08cf0d0zrBVWLBBHKRDLtKW0U9v2TpBIZLeYvGxGAekeAYn31Boi0RZRmMJvEfGtaeBOfxY2Qs
MH1g8jhHFq3PyaXmOMun3/3eIfSycF7hlB/TR5hPSoJTksdvYC6j9wGnlXOnzsxSEoHWXdOc97tl
mMdYinM9B+DncdY5WRVkvmEzKEiFQxNx9tcnuNG6NNuunoEKlx/ZulByyiMCnfdfm4vG5HEW0/4v
0VGFFXobtOBfc1ivkhpf7TwULyogNFDOTYpqcK/kn8okg0rP9/mRNAGC9QcvpLQkS5znen+HH8lR
NN2pE97dojSNdmPDUdPoaZlPele9n1GuL4jQT715WyiIgeYpIQV9S0O4zE6QMCvg2a6tjMvX/A39
ymoMMEIN1JFCqXcdnMoIQuTMuznjd0y1DjxcfZB3W5HviX7Ke8oAhBfuZ7HCbmwQ+qsfjrojwZod
q6dRnuqTa07kO72MvO11pvTqYGqGs9cKZ+jmlUv0LGH7YHuKe2FhXwWD9RR65wY2H1uMhMcx8J9S
FVV7smT/y06Bypo9warJdG8NuNBs9tmhji3Quq4ZcbAJdsrbhDPDKoBOZ7tjHb18iAIwODAdl6Vb
OFRnQUeF/lcqq6Xn/w9v4rdtYVZFDSRRCkznsQ9G6n389yvkJ4RWKXR1Cf+FfBjEMmLOzKQwUTqH
59CY7pDWFoh2WnNfRxsK5yEc+aIlzuPZbIiDCiE8K/3+WO3UKdT7iwciW3h24ylVJF7Sjm1iVBhL
2fEjVQc8CB5J7btpsj3SH7Qwb6OzI7ml27fTQsb59cRWsOnuIOOL2OGXI1jLWoVLayRjjFRrN4F7
dHBCvVPTrG15GbUlssBc9SDSg+Jwo1hR28Gq+Oso+lCmKcFRrKaN3Q2AIYoaSOEtrTwcWZ+EVh3V
F83almSTOSKY6p4m2RcCvkLjS+AurpaMOIxDoK/sxSwm78LA6sBgmc7qzdsgGKA91tBf9aEKm66c
Kis1u8fCA28oLVie04PGi+PThUp1ER3eJptsPXZJXW0RwTfBozGqCXy75jaUWNUAZJcEvt2CE3vj
cBe11+XI2KSIVubnUZ1LgCPeE5m8ulR04YZwA8atxvluW4zaA0n0opDX/Gmy5uKzb2zQUc8ES6Y4
eeXKh460Mwtvh7mclCwRpQm6FHO0jow79vEfC2FQjlEG+LZh1PVKow3JNeJb6YhgS+H/YIuJlgZs
h/8b6N5rX7zI132/WuqyBp35T9tk0kKHZWDb5306o3Ntnn6TxNgZqRWZXlj3ip8eVainQIewu5EM
Gn+8Nlniz6qnS83XLP86giNkObwWy8zJL0PWjsGGF2YelKDiPzZhtgGY1wrOBnW3cVXbmlWQt032
dAEbOswMY0lk3b9ldGfgUiiCPpxCnp4eBgrUgzJ1bnwDApx6BDU26up+/KKUvqHkEGD5gJMPUlFX
Cc0iWQGvGQgkekQMf9+zty1q/ORNMQwmHk4T8LjxDaxWRovrdMZWpWdBOzF1lbs0FWIKsFF3SpQb
wXEe3ZoN8MQ/yll/A2/wM9rZRwazXuq7kxSzuqtqwg/010714AId6UySvwI3RqVFwiKW5y6KsFrV
0rSgf/TVhKFHRS5LyaS2R5C1di2kIF8k2U0WhBXbimR7E6XrvQmGcpS/D/wULXurKVAV25R7gwTX
oxDxWLpW6dgnm28cIWKk65LeEyHkbg1Wi7aiXziizvhFdYav9rwSy9Yo79ZogtO9RlLeqqykuWPK
4+sNS3swv73go+hjTGid7t0N+OECKnmi2+T04XLLpTtheTadiF/cxgP3K/R2qKFmEQZFhf2ZKom8
Hz3PBngMuT5m3B2MtSOSh5G0Wo29blWJA8RtODK/Xbt2xZhALPdwV85rEYR9ueoe7vHWfB8X0Op4
/B90er2MJZ+ZhHivLm4KHQpRiBnk0aapSQbz+ode6Ueiiy/T7+7Q1+apX48Of1uAS1Y+WeF+s7RG
LFlu9ArUI1FmKz5Yz5zPAMF/QPm2YROiOQui75fgONO8Bc98IbTPt3lkD4+c5FXxvqRlOOt8Omit
65TXcI3uFhaIUU8ArtnH3LIHDJ9ZBif0o24WA3CZpNrNuOced3HRLvFd38NQeIW/PVPs2b80wk+V
R8b0QoWE2jRjNrMBx36tpTwDvspnn73cNdilIK+RIizoIDNwCxEMZnYS8s+62aBTLNd9eVthbq4q
vwTj99jOqi+KeFbTT5dGIgRDPL91a8e+0O/ux8xHim6IFLrQpTqGFixfs1zdyyevrzfd2+KmzMan
+EwWsKPa2OgDtRAkAcvXltvTLTPxxmg1kFCKPKMSPnpL9h9Rd8N4qTMpCcicP3nI/GaSZS6cFi4V
W6qkWf+Z5dVE5fBGW/IWy18cFmrro+lEXoVADsBxoMzfsWr2WG5u8DlC8hTZQcYy52kLGJdxiPcu
CYt0s4Cj1c33xHkxaf+wqYUwi6NZviFFP6hqygKu4EkmaPF9VRFo5sjNB536saUd4IvZzm2EDvp1
0/3sRdLIlyHbt1myZithhVRttjSjNi0hIEZ95BZKNcGbc9LaELy9rQze/ETjjPr1do76pXRVVuYq
d0Wlm0W1fKdoV+mWkMmqdZVU3qw/2/Tylz1yIIFfZsK6yGHDFaj5QvEW1BNFhNB1dJeuq7Yndyaz
51DqWCSLA8n0+mo8DnCnLG2vfA5QJp8rcQQuVGNKjv1IypyHgsxFEj9hHDU+88CPCPF8kGidWavu
o0KtD85IzNv1Wx7SLrRyqn4c91SrU5haCgdZcKT4bVLafw9YcH7T4T4cLoFjLFO6K5uwuc2er/Dq
KXoT76qAXTR0L9yfoA/r3zZvNVLn+TXmXvKfa2nr146815DJEjwEjM4H0W9bcWn9iBq+0zb1dClw
zu0Pn8065jg2bLCjLRmWGdrDGgN2YvuTypQmsyNPnQSg01d4dYUcvlNjBCATdAyWrewMs6qOSf18
31QsCtv447mWeYrY6/2xF5ZWpDFvu+js9m7+2Pk516AX5IXoNfg6w4igVLWWoCARrxpc0bTlhSmy
wh+YYULUbR1/Q3GKx+8rn3PogZcsS8eadpr4ttf4SA9p+7DdvJQf/Exo69Wm4X4OrJp+lY9ohF/0
cXHvlDFhkN9AeM1GyQhbFtiCHPonw0J2o1mB2UQW7s4PhkUZHdfcMDRaBlpWzn0OauyFaHSU6+VR
E4GgvGLy4KccsfLrjZSuIseg1BP52PfZBuPZ0DYNLhH3z6/aFilnhyuYgnLYmKW5IfgYO5LPk0iT
dp/n9bsYJTnJ5eGCGjjL4Sz5N+8eV2elFGW01FDeUp88XWrpShYKNeOJS2TJ30uqoiD6K32yjjAi
bIjaXMQTs9bMvXxU9qT/tcM0BgF5r80LKfE+YEJnndRWH+pf0eak2nK0myrFFrLV3bnbFaAHoIwf
2BMKOhJy9j00HhulGzTs7DB4f0AJW0dQbsZtV8cyDQKBIWGLHqvzv0BDfXE4sKIY9yqyHSaF//zV
zo7YDo26ERg1j3rODVs+O4ui+k32vkq4eiLj2mtTIiu2VIVRqIkzQ366wcFA/Tr/aCh5G10OUhwH
QKJliQ+U/vfOr/3hHEoQLYSt3iQwYNkA/ZnfrMwx+K88u3rBS78fAojbdjxZq7Uuxg97OXRiqS6G
dmsI/0SnFGVdhQ6U9SfriF9Lk6kd/FxpMbDK13o6eeNpXrNDHjFdL0itfbiyqJZR8RDMXtWOruMj
SvlkM4Ss0HRQgyOqdNIwWqyegh3lOVOnYrvKndVOXn1olBQpgM8BQSOqJA51453QnJXxtCbyx9lt
Is8+nKfDLOBXD7bOVrJ31soEZ65t39rHjIZv/tndhXzKVi46vGoRUzjKaDLN8mIuiVDXm2yEJncT
sXU4BbFxqRxJZ3nhwfgsueBXawfSZOHJGwaEe0WlifV/xLdSIvjowRIzmvygiWPmbD02dwgo9K9F
4vxfJlARoM39e5P8UhQa1cF4e5XGCjPaou0xdsONwBTaPIuqIbZ94SMnRIgvGitvtjOwelI49WrJ
UHLmEIeCZmWTDpEJozxkquCOtbK8y85MNr+E2kcpRX9OkWVXl+PuN7LJcfFSZUx85wj4jZW1bUzN
awg3LAka0enshwA+Eq4JC1/Qqri3aEzenTW47JHhvHWWAh7AaaVc+m2H8WSh7GyiKtKGVOS80rkx
5MOfSJw8Fw9jT6YgDUQ9j+UvrM24DLmKTeLtG02kXZTMEavx1VYnIg1MaNKo/rgiartzdXb7clRt
+n5lMJX1WeqOfY8H8rzFwZ4r7jk97nlogxMgCSZD+jCbzN7tGrzYrZ9cJCf1NbO9VV4YvgGEIcJu
tow5SNpb3rxjhvQbXuY4tzsMEiqz45wTz6vRaOxUuzKttGZ3rB9Ekmo6q7LcQ58o6bmBcBaQ7HoI
kt867b88u/NjLKbwho+RB83sfUo1r3Zcvpr78H50DHcG4zjl4HlkdRrL9er+U4zKWP46DuRsfbgp
BJe9Q70+ygOnOf/pXJldiYZr/pjVdXfDvc4aZZJadNhczfXxj4ZMA35qd30tNzlJWosIl0XHeMju
8K/w6nDz8Zgi2zXNTUyXju+0k8+Oy86YY3ZsJ5HNZpXAAgLxn6/7fJfXJDyyS3RbwsbTlUpGB0lp
etc2wZ8s56Y4CUZ0uusFAtT75zXxIgGRtVnkvc0eLUZD8+huzhq+2ogSw8jMXIAnbsPiZTHr643n
gl2/shUVZBKOHx4X3y0hTTYshCc71TQWZmOC9PbgKY7qDxjHmtF4BEOgWrQbY6fj23iIXQWYmwSH
ypjHHalnNuwXWvtDYbpvQle9CPFrnNd9RhPGuVSUB/+Txx3L4bE9Dh5OIMQlgpveUObcnpaWWMis
R8f/XRaAP6gCSMwaMqHfs62lma0DT9u1YhajXZHjM2fB5fOl3ziOpiZRyNq1lKWoxy5CTbzMT5yT
IMVVZEV6pjQCX3OGzpIzP9i2xoUUjkv47AmoZiygfUjqI9ILPaPZ/YovknKvLGXVz3oqcf94L4cR
sHbn10NbX+hyW3CYFA7U+4LJ3iZSlFgoDrFeQFzmUzsqY8xZcbJ5oXWXWRaWpr5a/OOI3kNBRnFO
UZDGWVth/hpb5YuaIU2Ht9SCd1ot+Lh73spv91XnHnpbVj0o25o+vNqN3zZXt539Gj3hyvYRrpQZ
S7J0QERc+L6tZe71MoaF5bTv7Ui7LqeHwHaA8lW/VbOhn9SCfTSzp/X90xVYBohvYGSAfdU59pHe
vXDBlrpWsDvkvXrHgkHjAIZ7+6R5c8//L6JDr3f2XFBAEAt9zD8B/mjpJZLnuOM6Tl3Qn6gP+IYx
VKH7VNyqrT6TS1vDDPfC3xT6WiEpc3le5V0N2CPa/9t/Ghq9FW3jCzK0Ds/bXjRkZyW9vDqZDWI6
dCcyU1L6FaJdJR1NARP/XmBTYrapUIragYp3JfKX3wkucRZ7Lnrjz4vWL0A4U3XsuZm4GvMW7FOo
67pqAzkVQnwGV6J42/elEwud5nSgGslKeDIATwek1YHjNVt2c9g1xFX6W6bAXlEeCi6klqJ5buVr
znHVR5oZFznDWqI9Oyn76TiJ2H6cktr0H+j+ohBRwtP0Q/Wwbw42gOex874BO8mRoozkuY6uvfWH
YGHCNm5f57KrJw6/AHCPbSyq8n5PSdbwbgkMQKK2ZGEgihgoLwmKTf35LCUzTkzEDyEAgywmvGxB
zixI+lOHDOfuHGuTaus55Fyg3XqCKOZch6056Iyky7bCrlWNSkv4oS7HNa0LOfkKBUYSwR+rPmZh
ju4oiAw10XWoUVmJlxv4h8dws9q73OagnwRpG7bHU5ZRgl4p6kbleoG1KrEi1+ix9eqnCvhuraMl
saJire0bBoood/Zj319zfGeYL2/FhiO2V6QQAjhcpdHJ3xrukYDZEpw1dd0YOOxmMhYk2nUeOcPx
laFFsD+2ukPV8n6wqMS7ujvbTHmFFgFlIp5+TSfYjFicyVkkvJJ9PFNk++cQnwZli0ad6GKJWAlw
rX879CGj9zQ6KpnTW2U4LjH/tdN6lSZ7CQXN3f6jTycWLZlIu9A9Ihemh49UYMm2w3SsiJoXrsE3
GBePvT16UNWWpAyVq/lJnrqoJLNjvNRoUGbdSZ28/mzjHeJR0bg6N6woZ3kVDK4Zylq7dM8Jbhxv
K+p50VvhQEBsCEucOSwEqovZQ1B7inm3UjnzNi6QVNDez/E38Exguzw8G99dzwYn0GxGrgwHCG4r
YEerGhqQVg7ExPZ45n0HeNVO46gEDl/WN4z0WcmHbfqCGe45rORdolv58KyCKDaj+/t9hMW6a5lR
D/RZPh0rZphADByLJvFIndqb7h/+vjKDiHys/D3MITM4sWFz/6RPRfO+S61gKzx01Pq4A8A+VXxw
kdA21VPdP51iR6RCJEsh8+Yh+AYBBxOCmEAazZ35I+PEwsv4m15FmLn46pXKFooJTa9iIibZQ9IT
tSSRanIcrdpVBWScZxoEJJPt3xn9pREqRmv04LhtHTC4IM4qS8LibPWgKFhSRBi2ULb0pqqQRmM8
FtRgirckRSUieL4BYKinjn3b63hLhcCf1R+9GM+9jp7whzb86CZRp7zgJ04wafRmgh23Tjk4N4bO
98bnGZcsM/vuSZQBkHF+IPRnZ8c+FK+dLDhInIR8ZlVBoYOwSVoSwgDHugvalpBHGteftHTOsDu/
w/43uKyMVJtUoGJH4ntHYW8nNnzGv0nidzzfTTvC3U5xE8kphDC2Vo7kBS2mB6bjWN05AR5C1D0h
b4XQBOkfMMw8MKefAa1zCLPYLA6VLJjWlUCH4je6RbIG/50kiXGNhIYGub0xfRObBwMamt1Cu8K+
deePB2d+w3A+n1bDHJN3cbBQ6IUqC4j6nXbNT8uyJEbButFczyQw+MxEmbnyrx2dVs8L6TRJoXZs
RTrjK3cgRGzMQcED25qEF+TcwzaKy+k25X8e08VOTwMQxu0PrJeFxS6cmCwIlCjZgR4hSlcc85wD
1f7q+FMjQc6rabbaQfEb0fKcev/2KfqPy7t1mfgYu8ADxyEu67znGGr/fwhS5CRT2kNWD9gKwmGy
97NjP55YjkhKa7G50YDfX0M9to9g4uF/7t0NoNqb1vNLFSjTTDsddCsQNZPKUEme1/hgg6XcgZcp
Xf4nhuMjNAu2XahE2p9Q24RcWh10u2FXulSJEQh8mjK5nPmzaJb7lwU5keAaS6TKWVI2eRWZaFHS
Wz0SrrInycufKAUoHP+YkRJwnhoHhQEbdS14IiEurbAsM0zhtus4bLcFjiHhHruSYAm9Jpudwn5i
I0pXLV6MHd4ozHBsVxamZ7IQ7N15BZagKkS1O2t83TO6Fd/pDZJJxSir+a2PdY/Fj8mgfvqUfWpP
Ih7NfDCQO2QiPGKA6ygoMNY/Tjl4UgjfBI0BV5NyKPc9fOMX+Xy4kDNJH+OWdViDnQBYvVAX8+YK
mjN7vwiKM1B2eKfRgyEkSfAEP77N/yh91etAhxaZIqTZZrYnsfvDQJ1RHMvu6MKAS8iqP+dqwP9d
FyMC9KRBYNtDRd+frSwT46Ji3YUZdXJ1P4iTEA8AYliQcOOv0+2shyBZrpgb3aOcCswp9PtyX78u
beYYpqyKJm4SYFWQHTRjmbWi0Xvw06gZWttdVJ9p9LLelT/1snPu3YbAWpRR8h8tF7KFjBnYeb5a
wwq7mSOJL0ZVmErAtw63lcnDTHjZ1ktoVCo1CzfLlXmdrzz1h15s1FwFkKeMJ8J96Qz3bPv6SUDU
e9cl3/Ydoni3zIanUtrQtw1tul/5U1s+Xygx6Mu+VTrWg3763ziuIneritMVC85HhyXxQTAz4tbT
PwjKsnLWoCo2K+8accMJvHFquxcwRhGNTaEr9lcATMY5/5yyBntHIDk3vPFP2IDtuO/fmf5z4I6o
RAGaqAu8kcV38xOqGv+1aukWACtZV4SfO3Q3Y4Fk30ULshYYoukxMfjCJ+6q/pw7E3FaxCrk09aK
wOW7BdAkYncew47HbS5a1jS0iZx5FBqM3MdqnYr2C/uH64wt0CCqUsWS1nVOtWlEx2ojT/B9R6TC
uDqCIwM0Tj2VN1VY2ZiYCH4PnCD8YX7lwrVE+TpV9xSc+OUIEfo0bWf+zJWARPe18GXipWFHPiif
sN0mUN8+HhCwzqjQrQT+ivjurHGPjmKDbSEYzL57ZyUNcXLWF33M5alBdaMqakd9rb38Yl0fwC+H
c6yjqv4vFlyrc/EcbG9uWX2Aw1I9qkQwXRCJjQn/RNal8BTU21Lp1mmFJuaTcoJisuzlgUtJCyGf
Ns7hcOGny4UWdVI+k9h9owYfT3iUJTPbqXcr9p9NJ4+loX7L6TQ/Dy14NcS5kZ0edn0V/eoOBI5F
62QxOdKmwaWgI8owG9QkWnQmLzsWSf3WaMJOwxX7Nni21wmAv24JtMCWqsI9UECRexIhv18wVdFs
iBKuudvFMrzAtNO8ffj23hMqc6EHN09/HtbgPeb3hf/4J3dpfsopflaZ1kNcf04AMLabHDctlekZ
1JkDcG3nhmnp0m9IGQrq3ixIP4saHuLXDiZeJHDx1nPi8YJP3IxS5H8H05ayoKhJ+UJ6X+yeOBmA
xN48y2uB/G3KjLj4yJ/m/OcY8nqtQ1hMOvADHUl/MGSzCBFhzi0ZWxFra0ofk6JW9QXuWmmG5h8G
tLO1uQcrGxQEnK2Cztm3FT+10HySM9WQ1956xQhCGgQwKkJNqgloohtxReMth7jomHUQ+6C0JsE0
ky4arjEBmZC4RAoPLMDNUQxCmFbm1jnCIylriEV2FXplr4xyLz6LCisw8Of4mD3SkXUafuZbFit9
GWesk/9qS29JD+sd7P0sqOSIh6oxBGrqyStziP+/9mkBO8IAFPSmpWWVDzytbmYHU7pzS9eiYVjW
e8O6PdyrpYEJmD+Fywc5vCsCks2etLkC7vuee/rxDjGiBQ7BqX1zBVTbH2QSww3t9mM9xPOcRJej
zjC0ipFzoiiKEoBVTiFT5DRbUSV8TdLfCZ3WzLq2pJ2uwjqTV8QdJkUCPj89j7XJm9yyJ51bbOGt
f7AX8fIidWw1Pd4Fu2k767mO71WcFl79RiOsubx6t0xv8rGfJxUYCijTT6NH7IAZnp67lY/wgln3
WqNXoWQihv5f1ywl9D+9Jd/7JvLXJrSNYM0TJgvR1mZooC34js5osFFmrl8GNwFyEUiyHecDF7vB
3qgMxmbz/lPkBFlvvzEhhFLCsDY9hqlbUf/IRvKFqB9T/xqR6EEdzltPq+xGXLUigIIpD9Wo7ysK
Vh5MMJMwarUlyH6be5Ins0bmjkMy3gm228dEXLtSID5KilZ8yJ15Hwd1Cletey+k4P3V2DtUuoaC
Aa9Yx+xGNTFE70lqF8ASVTHXxOBprT3myxTJbqNRR6nM1F8hzoNLtzIrT/lzaeLHF6GEXlYVFFfv
R+9X7vNxAbzldd4hUhs4rj8dEOrrepkQ1c5Fb3IfAwku7ykliNy9ocGL2M2y7PZ+B71/P/hCSzZK
z6zpmFckuFkTfl51kNcs9TkzWxsXYfn0i9MtAb+bxitBo7wGEUPnFadVLLfMAH9TmYk9E4zNEZI/
tHRf00RBKuc/VrDeiVyhdOaeznsFiZV7RC8JS6UayRqpvnqqQH+CZ1EV7+ufq3rnJ2AH0doHKfyI
HsKrPGMlOiSLlEfPiCOu28TF19h+TqB0qeuAgFd4tSJJbLH9Gk+nGy91piprZ2z3RjlHwUixB+3X
nWmoF/rIu0qTmLck5xJGc8UYxfxlMxE1eFBiGldkuYt0YipN5vfv1gkgsYuSEhCjeFA5kifKwYX6
VQ7GBHQwChDKNMdxtqXSjE27Win6LayTxggm4YgKgVDF4qIE6ZE/wxK56OcWoKWGYcimYkJ14HR4
4PocxpdYftixLWWHoI22c8jkoCmqrajfJ7DJj89d+as9j1UOnVsQR3W1Pg2rMCUxiPxIfgyZVicG
2uhALPt6eu4YqNDELJj+lFKpS/brN40F9+dCsasiA+o2PGkGhqX35AmTdpVsqMxEVnWxe/tUpfbl
nbxL/Nch+sUZc5ZQATvcFi9kyfnVzgd9979vGW7psnnZASPx2uWAZI9gJNQqmTpkaDAVe89o7Kn9
lNDLaq+OaBBy/JtNkWPb6fp5QgAa4/6E4R5u5D6jnDxO775y0zcMn17bDR27V0LOoExaml5I40oh
2jWlFvyDNRs1T4bsHD/J3bmZDqdb2Zc9GNo+S1I2tpbRcAGZ0pVQb5rT9v0E2wL5XP5O1PWPf+uR
AO5qKKXDMUTRkfLLPh4s79vXN0eQjIPqr7Y39zscj7/K6G2DdjlCl4m74cpxV7w7FZNaNZV8oqMK
SOWbogIJ96IMxMuUTPBON5T1VeTwV9rHgkV1JV4nom+5WRSpaNQI/6teTSvkq56Nf976aCYCyO4z
f/6L9ul/jmBeObXXb6KC0ZgEPlYySrzqRV4BFM2aGDyIP1q95zmBtPJ7jfx0FphCO/uSrvWxwKpy
Uh8Ma4juA7Eo/F9TkkD5i0JdhGHq++SUyvn98VZZYk7V4zV3oXpXUhJXK2zVP9s/0ru1h+9TLlE/
y80AVX3BB+hbQEXll0Yxtd+dI1ElEOZETQhEtw4D7ASJNdxrjZ9/5AB8OJ3vuWiIoD7p8qMpnSSN
cfy4nyBCrODnihZWP8yiIk9QOGAFIq4hYs7EWxdSfExRP8Q673zLNP5Iz8anffGIq5d25cEW+df+
G4PgiEIVzCKCozpnlyXKNA4Eupyio48UnTV97d+ED4lNSTX7q3VYgbWGNlv66HVieNRrTQsknxGu
SbPBzDjYRp/Sv814gdYyG+mvV2KLmKhjLcz0NhdknHT7tI30jCTfN46OPEEvkUFPh1Vq/WTOs9Hr
rJBoSohnKgGzkOh7lJq73uHtg693INnr4D7bTl+8FRnYayx/OZ1pKgVVP8mwr/2pCAxLYIrPYNGg
Ne24DurXnZ/5wpTIpmCNYfoUjuVuIxjXrj/IN/J+SGApZdxxvxeXJkSwvt8Bf15kTkvEOCt6Feyg
xpJ6bT5uAQfqXVGFv3zrN+0nUV0H5DhrrYW6av7DG49BrAkK595wEilWWLVOzTi9KtueeopIOz1u
QJKYHzt5EYDguHwGM29Va/JQwgu5rtHFgTQMP1agEPPjWPsFfFMzPzCwaDhi5BDIwroqLknRx40u
yCglHfl/+yq+OzLWft2jkEoSCaRV6zUDs4O7Uj8ZCQj0nD740miSuiIExPofOTuZPLK3Evczsstx
EeWjD/u6BI/j+XiQMfwYcp1R9d8whaHX832WyVWLNMG0UFWiW2dj4sAlJPecG2lhxk4dXQ7xf8pe
M+PQCh46E7tT0Zniuu4rue9M2MB1zcLQPUifatPYsLnz8qo6YVBpLzKtZRa0RpR2Voe7W3tRnmxn
KE5xf+qIYKBBiDqgDHQHZCYVowcrUYcyxVNjb2jPqrGBEPYQ232E8r26v0lkGPChZb6caSOxpnlS
oqnWU+K0dGYhCdJptEkI2En2rdfLPH8CNpBL8Sf4IDE+7J4xfM2x0NlmJRRaL3J+vmjMuISHmqDb
dJEQ4LRnXAR+eXEZuXUYBqIKmKT14QSrPjv2IePcMAQBqw6iS+tlt/UpARud+lwI1xFntQ56d65n
+W4qZCef2vMAxNShidYK3YWwUliTFdDIi9yoi2U4mpLOdmUQjed45KDrkpMfWB2GeAbTYF2y4bS5
YLkERXd5cGHBp3sUZ7YpZNVgEqAUzeQsb+0vMU/Hio1OI00AAQxOffR7KzbMlaRtF/jIZtx8ad1H
mKc6P7raXkn0Vt6QH/x0McROxyHXYc1tDsZdl1Cm8PTmes6ZDM/4q5Ahw9viIDYh4bSnGriiAKNV
zLdOnmpCm1XwBIQDsjmZrDyDS0y287Ou9wijM0c+0ep0qkkSvTDIMjLAQQmXiB0g/tsxLrxrnPJv
4N1sfHc3MhQxIdVkgStEoUW47saODbIU7434fa0aBS1cjkOxqaQNDCmzYKrfNSdENxt8rgNhF0Il
bBTP1Nd1wCdkZMx2eNnkjjzdIHBC1q4XMttrGckTBgAMVXsWKSb3ijrzavneePdIHmdJq9rPqnaO
JfSUMMWu17NNx1d6nescyMu7AsDVa5H0gb/STDn1YlKVgQbjwFZH5NyncUHkhyFR7MeKfXdck57K
QXQAx3c587zpD0VQscyAlqsj5qiSq50/XbE/uxz6W1RHEam1Wz2SBY0c7N6fONr8E/XXCAh5b6zm
UqbvO6uu3ggqtz2z0yCyHiiyu7eOGmYPEYgG2Vs7/Cwu1ydiiNSXUPNOvYDwpewrGI/O9txuY7Ld
DHBVg2DWovFYGVgf24+MeSOE3BzMI6yl2xjQS2mepl3UXUF/z5/78Z3lLeYgn5I4MEUDJN1m//B7
5SithvOZKItXD7yhrtCF0yrnOT1/38oxeqiZ2kkGi7g5Al6QKhCiJDuDnlipg7Ih0xmBoCLYZJFy
0w3zqRjAQEdAdhgJqwp+ntRYq5Tc3mI7XYSj0h87K85jwzmGzDuttMi59gbAj3ppobkUP3jjChQV
QzoV1npUz1DeD1AmnGaU3j52GsyjKZvUj/eLb4xF68rBd0Tre2rDIelgMrOcY3aAtKCWLbH8LEKy
v7Qzik6UaB4D5HKLBsICF4upy0jtAPwr/JdXdkUyUxv/n0+icYinI4fwzb5teV9PjdnmrRMUGpYs
jrq6MWwLHpsbNqefJGijlidLxSfHZg+UwLEw2dR0Db3+cokA8Nki3Hy8k6FwwAMJ1qd2tpCnYW98
33DM04pj4KEOyxeHmUfQMa+q3KTKS/5sPIjlSpvndmKTC/YP3Y0M5vHbbNM9YfPEajgbtxI738/y
B6fRLhs/OAJEgKNZYUkZXJF2hywvN38hQ3+QVL+RqQM/TA+3S/4lFjLwDp5MJnyxf6PaHNuDEUA2
NoFrScbeVrjuy9SGmZWpERkaMP1yKgjZPH0drsxOI1e6IhrANFelwJFfDOJrdVqvo4xBDgOMsNFd
CNyVZSRu/bdTjZ8v6Im6Osqd1nSeORKr6Enid31hasKfUAqyMUY6mSThfeQg+cO2nIPnHW7QHPjm
6mmE8ZEt1nF8sTraZ3vQO0urhmVjX8trFgp9q8LSPSyaM7vIGPiO66O21VGrR2qOIDPNnv9DFUpJ
WiLQzgjDq+a3RhmrGGrm9CKe9lHnJKdX9AXGtOmKG6exZWkRBecUUuciRJx5q5WtA7YmaFxA3H3g
AiG9SS8uqFr0WmkousZKAWeeawQLt37PVl3801bP6IEe7gNc61++LcoS0TW9IHgCoJybnuL4xVcb
0iTzjUUSwhYOaUB6bFkb0iRYLYHH1MMr2rKNcDtDmdv+9zkbkr3oxPJIxh9v3C/aCgBDUJs3Ewi2
MEIPHa8nts1uRmWVjptwC+0kleh7B8d+/+zGqMlrCZNUUGg3UzEHCPzjTFu/N1qzge3J8Z4U2Pk1
KDHsX9AUjc0nYRNjxIdFN1mho47PGbtr3Jt8BVJv+h952f+dq1waSInMdsTjLr3DdgCY/HX8cFwE
vpCuZ+0ddV47SkDGtGV8hKLJSl78ZMg6YceDed5xqNtXiS273np4/u5/zvAeIDMrH//TKBPcX7Yk
hD/NV2yHNGEXkSFd30xfBQPbwSHN896IW+NfdxlglrCGchl6W6kFAnagB4Ujd3TybsInGe86c/PQ
xr9ZQFZ6s/MuhCkrMilzJl1krFOxTpCMk2SGUXdvne07FPqQTkK9A2g49ICE8kVBC1fWJgnPqdMe
vV13pcRAxqBSjejGNr5rHqpUMxCOAsbrwj+ke45MYTnCLBkpCXy7Zp3catMU6miJvhslrAksUGYw
RvUmcxBK/ayxETKtxADCwIsDTAQoLIsa4ousyp4qKEvFZA3wNtSaO5DQyeT7MH6eOkVnq1bvvYPo
1BOkVwK3cV+yy3E75LschINgsR84Rw3DrB9w1yja3utmGtm16dxcxwO1jRIqrjBbDeSka/xkO8GN
lVYIS5RZaLSuwoHvNnDMG0WXoVbeYQcgIsxCxt8KDfY648600SGh99+h6CIoZ1yJbjotdGbXZKPa
Q67bq4D5LX6LBFsR4S34731Xt3M2KxKugvltdpotPGJlhBBDY6OIuUl05jnDYahD9zIr0oL5RWVr
jjH8FpiwInlmPCf0bgi0avp8sK6ZUEWQ6V05vAPyTCZcVPbx9lpIdhN/zHWdD5vKlwVo7lN94lvn
ziLpj5r28ClI0K+VMEh9i4KL2kczW3gTRSaHtvR8DIPmrFoitLxMw1emi0Mnso1O3mYUkvb3/Noa
sqH7fQ6YRXX1AnlS7T88BogFpC+QxkI/w+VFbw7WYFyd1GzWRS+rXW0FAap/SYsITrj/MQ/pc2td
v9ls6RRtG4xBgUuEDnYtMRcay4IXdd7+OQ3F1A08T6P0oPgsspA+n7PUnmP6EkHM7dMenMEmGql8
Ktfw3glWImAk3nUcexblJ6N7YVQHvR9C3e7d8ODFNFiKHmQDbJv5SuUmHKoBZUsqyTCgWQzfKQOt
T3iGqMoKUW3pPZnE0dbfSYV3eHodrL/7yil7THMbZxsPkwuTFFdTwxRuLgxw7MCdM9UGICMZ8ZEK
55tnliTWBLoUr503Vjr8pvwikpCLEnRFTAWtBlsGjGPnd/Bc4Z8oXJ/czVB112Jr9xErq/HjlNhR
J0FUSvoavGCtBNuxGRq7rlemFdMbAalOuENlrJlaHWMiQ8aXJUQxS6EeRch/4pjHHogpNAPwxU6+
M7KhfkAkBVZiFdqBsZDPvBl6cWQ4XhlzSxlbb2/7E6tIYehZob6hqKQ4nEXV9DUxh7fM1lIO1jdo
1gI0iBMlJj+5Zz+nrESyDQ8aBXeb98o02HGPOHag56O9gWQQL8tXH03A3Vfpe8ig6Q2YquOhb3zS
/HGdPJbIY9d2qwXbbdOhorXaTEQEcT3uzLq6c5EFKwFne7LhEERvFEF0nmHAZGev8ziiSKVwBHoV
4AypydYgXaHFw6/aNHQtDl45nyu/QHahD+3fw2iiTCUya9sMahlpfXmxA+MyWdNIqqgOWTPOmf2o
CQCm9PgHLghArYRDVlNDTCO+RIprkWH+Vy5DUx5QPPylY6IbTiVjOXU2dcHF2k2im06kyIOSDexV
XzuR01zd9v7uGK7nSN998RcBPqqfMycAuLi+VCGxVBozdSLByPIV5M/c/K4o4DQf6Xy7LwOuhHDP
svO2UKRkqAJVg5SpB+woMjM0Nu7ts+WO+dS3vvAnv+03hS5fdmasp8k7DufdGiy+oOXK+NdsKrTo
w06VRjr/iHhV3ih6Y06zg7vIArpEUufFijlITflZMxY64Ya8tW7LGeb8CtPDnl9fo7OekupBUhNx
VdTqginwbyiQ+zbF/y6l1E4m9jWEGl6eEXOxqz5Xka9agFjrYDoSE4MhtMBiuec6+iJ8uwq/fcN0
fYOpo+hCaRdIiPwRr41aVFRLIqGf9O6Kk7yDJ7qs8A5+djy3K/eAlmebODmJnbHUB1ZPq8V/YUEf
G/VrgxFJKWzU4p3xPc/ZTVCfh7csxvLx72/1e36fCqwTtQXuTn3+dgnuSqwUJ9MtXmctjIxjkC3s
LXp4IluflorNKtPBhkDoBsbs5FIji/NuUl7/fWqiyBOrfArJIrBE4vT9Mc7MzPak2x8oZ7LPg91U
iE997UZQZhDlF1YgDb8FF+z7a64f3zzkcJaHGuIrg18aSMdjr31V7DDgfPLeYtK8YwfmtONw/CPE
3ZaV9U+QN+x7FW5PMng0eMvL0AI07JtaxwHraEGJVUHcaWiDnamlx8Wva3RAexVelJLWTvlXwcBJ
svuGBSSE+xJU57DVVZ/3YkuFPX8UYSeDIXUed89WLaKRqK+4vDuf/aNjxV6muzaAHv1FtNQ4070e
J84V1YI/PiuwhK5mg6ev45mSK1y3gObXASQCAVz9mKh9CBc3v95sBgcrMehO6ZVGkxU1m97SmLlr
55bjF8AjKUNH6s5zgyh8fZJlCxp5HAB20q1GLLkdDMvMKkfWoe5tdp38Jz7jmkDvQ/1dE7ZEL+/Z
XsG4JrEItUoECIRRzAu8Xj620dFbYZmMPsoDlLZCqaxyaglM3cen+Pz2A6VHPP1IanHaJe0WICmR
vvaOfNGhIPFHL7rdOzeuVyJK/MOVC3KireayEXRdQgk6mr/Nx6jgpFJMwuQ/4y49DDRSfWZZLZpZ
X5ks/eay91+2V7jSKkwzH3qScaZZfsRxa5rMcoBkzLQmLCrU2dyUJtqkxXxzQPju3aDYbH95oI4l
WviOmVx2OYuo3RXWGFrIrp9zgAZo5NZmzomyYlDD/1VznzFgJgTQVuCgpCVLZOmMRzpIddM+/sPv
G7n9bOiDMhaIbRo8vIxWGqLaw8v6p+zJn/iJKFwu+tE61MuYcv1w1OotPKsds6Wd3E0TX1JYBtMQ
oOfJGYF6Yee27n1BHJNE3YyeWck91xYuurviQVkQtS60Oz0jFgf2Dtyh40YQFwr62gzqe11YnzGn
joBzsSaxtd5ye6+JN0nIzoD8GmpEw4pgIKmaS3aWyfyszghEOMPVT7NorQlhBGUFkSDVuOiJFO/v
GY584Ue/3GKgEZWntreZAxlc/gGX4CD0TJXfRoLSbq2J1flCOLBH+p/DMHMnCJ34rxwNCjkw34qM
IyeNkApefQ91A4mRJRZDw/xsiP4oav8+27u0Rmv6q6lRzfWFdTJrPJQIkoZwntavtfXuehUh0rP9
up72Yu//i6OTkg0e+Kq+Db3M+ggtfW3O2oIOxsdU/0UTbzTKDKJh/I53NplqTHzFMdPvckZjC5Ry
zQl61oZQYlbz+4vq17S5Atxx2ruBmSYvfBH5kEqDUdmm7q4z/bPPXmYAjDCSEHkT/9N2U/C1jVc3
zBo5dc/5POQe5iuNhOBLNjfa+95UjBdtImuLzkA4dTphGifDlQcPeZfNmIg0GnBtSQsYGUjZkivg
P3cju4blEW0ZuJBnIJ0Pif5jfu4KmrfF9La6IesyDhiWLXpbZuEcE8oJGc27eXMjSgIFwaAIE0cS
rzNM5Vs8LLfxLZjBzRyGIenhluyFnq38zGXYBzh6JAi9NR7Psg30jE3xD085nBSMgRlkQjW6RXMb
jvZv7juhTeJih2jaKuaM1Vy+WlKSB5dw369yoi+aFNITctFV4Q64zHNSqHbh+xsxqVujcbCTK5I9
taUOIt42CKw2cbUD597WZRGBiXQL13BTtW2IWEYCkGqywTz0HsrPaVwF4Z20uHYFYImCkE4Z8fO0
B6yoQZkmQ4YvX1OzgwH6BeFx4xXgT27fQLVDor4+HNg4Et4ye613r3TVIwO9s1necEYpuOU+KGMk
RaZflIXYI4r0pM1Nj9WoYM/pG6bvwvmR1JF76a+iOsEPojAguxs72t/uCKpqZWphnkBcYouRe9lW
jRB7GWPKx2Iw0BYEKT8zTfBwVVB8HWTWTKE1jguTG8J5FXL8AiUtytmsVS/A/RO867J1Bq8JdZbX
C89wr/gcJ4VayGVjUHJy6SlRLHw5ix5xqa8nxpOqu4d5X0W/lrpOJUACfDooXDb7ztqWBNYcynsX
YZK2482FyTwvtxWOHqjhL42tF+mh4hywld0lISj8jD2SWLUR4VK2XBiUw2iPp6LPIH4pKBFcYoch
abP3u5Hjtr/zHF2gDageP90/mX4X379+7pg2aD6TQ3HIs6Fq7pPD/Qe42wKxscfbQB8dbLhUdz3y
+7MiTBTfcIpbslvf5DuOukKY6KEknuxEqhjqv7KTvUGtkT6aZA+/7iP7z2pKD6epnI2C44hB2fV+
VFKi5N1xdB2k3cydAtmF29fmu8LOXzclWXlyLcMqkqut2k0uCUwTBUObGM6PEDphdx0eaHMJRvW1
6foRQY2FGZF1RBRaKDXZKo7lQeO+czomhS5OOGCTeVAEJEV5D2OlPtWOfoGHfNISldQmk87IAjx4
E2n7e4GlxWeyb1H4pyyqdrrqYgFxuG1s0wTpCVMHKXTdVIDGlTOTP5aHWRN3ar2UTUNO+GYCnmPe
zhc+nJk/xIH3Owt1bNDjvcvwz97UOK9R2aLvRxNHvh3FWMhXF+HxeinwT29ZV7aRAZO6+CCXx96Q
yr4yU+eIXDXx/AatC6oXSolhVWcEk5E/ZhZoZq4YoQAa15z+/lYFcs0ITNCpzMEJcRRm3tFk3k6R
tJ1FQALXO72aKOG8KE1/EiVe1qSXFMnrQo/vmk+mfkLY53GDod1qJ+Y096AMXSDWgPelXaSHdf4e
Zv3pXXmaJv48tJYxXdwdBFT0d5tbBAkLu2hDWnnWIb5+jeZgtMwNs5Wg/+E2zGOwPDwO/RH4ympa
Mwar+Mbfu10VbQL9BT38PcnYH7Z3LnwS5MIeyk036Zbu3aSho8+ErbF+xt27uB2f7imFuJI/DaqT
J5UmeJPerulJZYUEo8VpbXVibuJ2P5YW3npOKc9pkQ0FoIylNEOvKI2LKumvjeZVwSqFSaISF2h4
at7OzJVZUu8RiBAClB8Jl60y9trEPYtLRvZIcHLODIKRvYDmMXKTwMzdERBfpHcoXuKBHXDg70zm
DX81tZBOKW+xPdnU7TFL2sXn/3QkCNSq3El76hWHp0wnKqIinXWVbUHY+z9dKH6SBIkcl+rkTrVL
QQO0kY1EZ5TYK63lC9moHi3Q205JfRuGzVhc3APj2p1ZT2Zf9vIPL1NrVv4mMhb3GCJ2iCJ53CZs
WlTj54iKq1mZ2Uh4fppVSmBxZZnUWzxCORTLYZhl80RSks6jtyvu3uTZPfnlQNlm99F7ATSWoG7L
q8pPuh5JhGfGXW+P8Qs5MIhRge/Jnva+0vLR2MpfipvTnpoFV6fKm64dSVR89i3cjk6GPVQyP/Om
DANYkDFr2mtUQ19WXxK8s2ubEJUGA/ib95c+femB7do9/k6lU44k7J+hzJVJGDR8r6GAcVKvICTj
kY6rvX+vynah4yXuHMdjrFcNH9vlvj0WO476RQtTvw8/FizLJSfsZjHJmndWyWDtoVVuhV7jXBXV
YrAL+ErTkaQHmhROU6JQhc+XPwZ+PU8Fal2Y1nHoo2TaYAXNQ8UsZMaJmin641AiZQZk55zwSG+E
wXOuH9pO+3uOKrC98z+gZHmYvh7BjJBvteMsPNcF8TUKaiTABZMRqXq7si6ttcH8wfCyyKr/o17g
iA+NqyDhEGbF/uuPHwbk7pVn4qSQcgQMZkQ6AsPxuuDT+JXrkNkmtSr9Aqk4ZiCrEO+YgNs16Pnj
KZOU4IefLoosrykQE1L1pI6fezGtJlopAPEiTBS8yNVUPRNQlX4LWR0DxG+qj4H9fYfZ2+/SEY+q
ewZQPM5d1kE5ckWngg6NYpxOoq4xQHoIssi8X0dw9rHfEsmqREqZgo19y0cZ0HuPMAdH4z2i34EZ
9v/pCEE8ebDPl+mPoQLE1OYPqifv6KMLk8PIsEatDAwC0b8FNUg9O+A34OpEe+JObu1UUlV2b5j3
mQxcHTWs/ORmHcqPBNwMgA2/yz71ZlR2SislFZqUQY6jV3uQ7xHWpqJMSqUUeYtYELaeTCfIB6ZK
DfhRGm9+TBcuFFcYOkoKPfFJdgyYvEHfrUHubigHu77vlG+VcJkcrup+Qc3Uz/KXs87bd3QeRp6k
Dt5NaobYgoVqlv906LrWf3mevt173bjgkT08o/+DD64qBG3NiuLju2sdhi7hl9royt31dOEqp8Yc
XCM6K3OnsoO3reYmSL8yrrvoQ3jnGu24gpOztP5CGO+Vm8ScJasGQsemPQtnBUXUC87pAHyPBKqN
b5alErGIccbrbN/0N0p8l0CpitM0Y/XckyPbkpQVJDXqo1VGzDy8jOVi0qUnxNyc8eNxFjtio0Z5
GT9eIpiXyRJTzz2RTmCNPvjIXjbscJLCTMpfdNhqVSkkJjGQ9edBOvJi00t16o/nJPwVdI+HOARX
PACECw7gvYz4rvR0JuiO1K2TlRcGWvVogAkz9TDodQCO0jjouOC+5S37XW8X4mG4sQKCNSRvtr62
VH5nfJ5/pjzE5bS8fwpbgD13AO420ME/X+cxMnoAVpz8kw2RNmNNtfZHIOoq1YKTwF2cMl/Tc6MI
3WmEDFsI7SQjf8wdKFl3MdfwBO/KMV/+Ry52fvHlPtlZ5HJlna+RG33/vUpptHp2W7qZSEPn8qoI
+R2asfTGKyjkfIp6UBJYGKPcupI/b4u6q7RXO3L8k3Z0HSwcNs405xyeyv4mlevG8RjRirWGnIBz
TrQnuPqFAnfPVOzwbjWjQPrZZe2G2axgWZsVQ3El7e7QP9fVEpRF4kLBpYLxQcOyWQVTWmw8QCk8
ahB3ixNbTA1Li4/ZY/bMpoZwdwnT89TrSj8fdoMWPL0rsgXwJzsQnOIQ8NO09OhHpoGY+HjnIHhN
T0X4MWJpk8G12RgRTcuP3LvMCT76n/Rvp0qShqpXTlac9jWe8KlLGjStPz0RRZBfWvfgYNWrnC3o
IBxwZzlQr6LYLsowAQDtWA5eVYyV5sUEQzm6UFvoL2hWJxm7ib8Zqdu5IHdm+Gx5Vo5qbCGMggs+
SKxgW4Qka/nJ+BV2ZEwWstH2GXZktkE7iGeam+MjkqHSf1acsjJbDOMK+qdTEn0grRYIAgRrL28x
LAUmzO4IBDqxxlLW/ZsWyCR0nZcwxu6c37VIhxHpLbbcWGH3dumKMSDFIo7YGiW4/m+1C51lcSap
hu4h9Ypv3Zn5FyBl4gSs+4E/SSUWKihmKKQ1uMSp7JNuay4OH5S1I/+7dPkDLTV0I73oM81Fwg2t
K9ZtERBl0b3Jeta/7rvQhVxIHInSIUjze2YvGGk9MtU5AYOjgQlHx1jzc/ePIvuEt8U/aQi8f5/b
Ui7b9Nd1lzU47c0VKUbCMJ3cglnlpIXf6vvO0wJ+XoNHAFHbwPDZruS8R7z626PdgpK0WyyxBL1i
hvl+dGplypm7IGEdSTLTVXl4lVT788ATUhblQjh6uPkZEda+G2ExVoRxZdMZ+gyd+GwQf3xl5t89
qKICZJY5x0RE8qlFjsWQRs1kzkBejPaAPc7FgTEXlI6LFHLICanizyqFwrPqAJS0jBE2Xm3mIw2U
e/YPG7VakHJ3LJ0Ze18+sgXVQQ5K5fcSHEm0le8ZTd/KGfsryH4p68DilLdObn72r3zJDSs0dLs/
aPHJrCVvMlOyoAdwg8sGb/YAHtjxlBjQ67rsiBcUI2zFYDHyWJvwtq1X0kGEM4sHN+bzFwrp2VR0
QaoZk98k2L/ySvENIOMlWWu0XipP299M8YGfeyW1sdk1+gaOI6stDngcGKKSCuxkIkfp3qKpglla
3yFkhOhkfbGb7HhiGfqVDgv+Km2zykWV49SDN/w7XCFpCmNGvsuHaM39E5nF3EcRsqjNZjIgrVkA
3DysT8FKRCQXdIxdrE4f3hdmpWaXPqR8voBbThVsJsLUFIS+T91GS+quubE3+ikinggF+IRkHdxZ
xkCW7BsDJfipS4cQ0H+O4tEWxj6wxrwLdeExVbsAy8IrFsAH/6MrGjbM8VnB8f2u6fp5/bhgZtd1
Ro17+qZUzG1tF/CjtfMPc8vRC4MjKTg/SWZHPNkaZXW83ulYnmQqqo6wVUozHSoGr9HM2XY6BNQG
SY2ABl96iogbHsM3+C42mi5DNl3Tyb/EChNDIAUv2SWSmm3tSYCvCWmDzKV82RSyyBfwRC1cv+PA
JNTKjY0aARPOW/zrjAIVOSU1lqCik4UcKM5aDzBXLFhKx/mH9YWWtNZB08WQkMPspMy57P+CDT9L
Lg4el6XnBeRlArGc2+ZozaNZOqueer5oK0oiA983qFLdakjbzPFxNv+xOPV9fijX7o4BZtSiXH1R
UVsRqkPUmoGnUStedFDW/JzkAyftStuaWZMtXIdD6flsRRVHN1/SZsNYtPABxRgwM2MVoNd9MUuJ
MYtIntZ0Bb24fripyITkmxwOE/S509nhN7bdl4iUu4sy0Tc39qze208vhdN7rirC9cEaWajsl5no
lINTK893p69DMAj4u27yJ2j8tfzkmo7u7KVL0vRUaw6GWybGEFtFiugNCjZ2ZrB6iIPV+nM+wOKH
8cJovTyyEYqfDdZuEo6iWdKdwd2cMSBahNxrCfX3aJHihRyyMakyFjp7uDD9H3AOhkc1LFzHjVO+
0HEeMBq39k8oxQS52IxhiX8/W8ZGSKbO8MleP9a6sbGQeU7/dhC27EeBCEL3WGBYfxAf8uSBwXZZ
o6tw4tS6RQT23rVEVH6cSp8iWLAgFO52Z9TJskV8pm2u4PodVxbZ2hVNmiNrT4XiZacdmYxM39Ui
fX/kMzXhmXq4VGSpCiFYeUsNARZx5WtWAs3KSiz1Cozb6jxF1KREI5f3A5MhBfAOkb38XUwz9CPL
e1mcnipqPqrbwqYOtL0sReO1RtfvrUUHptnAot1xRTavi3mOcqmoJ5AeYEm4xdQqZSmANk/cVL7S
6Meqoy3V6c6mQs1Os2jK5V1dLzBByv6jYwlCb+0aYbO1cXuw4W8sh5FZCDEZlTIYBHbimz2tXNg4
9XQiHuwP43O3+K4Vn/0keHoKxSobkoK9a99AvMQ7xxnDW64XxxPRFwCseGMUus0K7yE4SDMu34Eq
M7IRIHyLTWgt1TciEDuv7tIc/HlAQn5NZQcl3pPCCQEwhE43TpRz7Vy7G3RxfBsl1MFFKMIFemYR
cc0aGBV77naQzFhkoVT5nku7tX5IkNEQ+C6DEk5K/3QrGX9LKU5ti9aOZ9mgAijAFswvFMXQ7vf7
n3zBaDQrc3oqh4LIk+rxNX9QjJ27e7xd4aJ+4UYjM4nODzauCYe9FZNL3hOLJyR2RevdQLJeVLwJ
GWDGSKIXuU4YYa6FmLKX/IbBQi8t67iUCmNO9VEF6NUHuzA9p/PUWmE6NKxaY9yEjDknoQ8T4Xo4
LzIepstiNdYmnqpy+EVP6aI1hnribLWhZKoHcVcY5y+BspJDa/KtnKp5iNYccx6ckBIChDfmLg1s
o9uYG0ku28crkVwo0zmXLUi18nKLlYhEJ1XSVm4UwSOr14S1UrudloqtoXkvDsSG/QzBUTl8QTvO
+zCkoOrzvE409aszJvHZSAfbyHcjYRcolBysTts2bsoxZJRioDiWyQ1DuP2S5t7CIyuhGQmzUY94
ehhD97ZQF+TcGMHi16LL7gqO3H4JCNEEORdeIzPonAa+crmERLOEF3VoTuhgWvITLnQJwmibNjuP
8NtqXhk8GgdNxWyjx5WQYLXFS4GAUZvwTgHp6XsP1nfIofHPno+HiLv5B0vnfrPNSwaXl8h1AnYA
0U6X1SwwVooB/ZtDGEIDqlbLVfdJkMzcc3t6W06duiP9+7hiiOC4UvH/CA+2XhF+Vgs3M853ZwPv
z46BM19sotFc5+Vk+BOwodWukkNZPdmjYbhIbheF4cG2IEPDji3C6BoSXue+j1uBcUDs343nRCEQ
MRNORm+iG0nmO8L6hrT1EGYnXJy0xrkFEHiCJmH1v8ZX++t9V7ci0ucrSLmnbNE2AwULNhaoJCwz
UxdMWz1MYAjSTp6wraLBb+KTZaNimXyxVA4rpSiNSCVDNr7bzA+ckUADBwXe00ZCD+m+33NIcq2F
N5aGnHBJ65LsW5nXghCOTfJD2KwO0NmcZOy5iCz3x3aEzjelEt5Vlx8zh2K53wOaAAgFvgKiVZq/
FoFymLl9b24lLR4mkzfYsNF0SKxlEQPyemweuky3ymHVwvDyjVU/zf34YmR2B1nBcIzv8bocnvn8
aoozo2N7CFp4krEy3pfkwmawPntA9g+VTysy+NA2nvl4aMTs0D/6oUJcsmbqr97cy3PDExjpDZ9q
rQOF8bjNqAqHuRhjY3IqNeXXq+19gQJwqEaZ/adVbKYqxTwqaDaf8p5c4zizYJN3Srwiuh+fmOnA
D6mzsx2ACPgek9siQGhwN75Y/Ij3/SIX1yqZzIw5JKj8xi7KLnk7OvXFWZrPTzuYkiSIqJkZdNhR
ZX8WhCetSWRBmtyAeSQ8rEfgiJWpHBh6uit21WWLJdKjwGtXloj97vaN1+M0/YGODYdnvD7j8NqO
DHYWZ5K5hwdCYrQQc+aJmq0AEw1Q2BkRPAXYCqvNEKWEdncVVWXKa7H1X6nNzliQIH2k5iw/aDDR
Hx7NsG1R7VN6A9ZttJJVpzFiXNZEG8tMtdGwZeB/zEBozilQrhV04uAk5tQ3cIIT3H4Ddz3sKnk9
TPPZBn24uFaC+fAitZnlyMbTiALiUmmuD0LPR2UGNCdaZpriARhlZOxnJ2+rtRCLA7Dc3Y9RIc+c
/suFeltC7/Yis2zm6prG85CNlXCNZl/0G9JpzZ7BVYKhka8NnRUETMnctLFHMQKMpYU9uGDFrr1C
O7G38CK0LwlDGjxkOKzKQaWVhCEsLEdpNbtc3Tk3rSH2XtY0WZ5dHVh4pRcElOdsqJX2Ag88vj80
6v2r3+2nnLx1/bgsOEWoUjjmLsM3jFA4zQziFcmAQM8rsYZxKnc6KJHz4oXo7NH8pSE+53xKA0zG
+ltmIv7wHrMRQKJJizLo/27Q0rT46NpQz4hw6byO9M82w0dIXNdqleNAKw9hvPWxKG/cdUbauAGM
ygyqEjDDVZFWaA2Kkm5FalcRylMaRO4lxQNzLbMlFAqdjSAKt3V1y+RazxNlL/lKW0GI8Tikzwhl
oxyz7E3q2nai66QnJAZvwwUuxCYP+QL3bNvegsY5H31zoIX6k4zRuhdLWvE662eTfk9tSgxUx3zF
S42qTl8gUM4KHW8NAYuwx3/f50AxHGIkFd305lXR57izEfMC1aV/9+e3GT7LQvTRN5Lzvdgv1gWY
RBuN+jNP+YP2Ez0NP8bpw6xt0mrKRmjUaEkFAFXdEj6M+5GJykjd0EzmrRFuGh3Oyz5fCWoVpCXR
VADjDVPB9Rh3qRu/Vw2G0LCugaebdZQkuOruqsAsmTSr8+D6CMi8Uy3QMV3/yEx9Lch/+6YVJza3
7Z2oPCQY5AB33N11aXrisy4Je1FUwom/YjcqOuvbsUIXJc9eJhMAUPyfjh4OxZcpLli9bABLwc/L
7jNL1ovrZeWOB/swAErfiHt6fUQFSDEk/XXAubD3AUNoDT5W3sFSgQFicvQKZwcuMyX+6F7VWooG
67w7tmeO95iXA/6AzszZqvU/m0iZB3gsJ1e1f7Z/1J680XN4x5q+W95jy7Uqpp+tsOfX4aoq4KVK
0aD/4I9SSF5F3lWWVk7hg0WjzWWVXUnCTkcGlPuz9cAgTFG/jIlB+2TYUFJR688qOCwVH/CbwOv/
2hf3l7Z7RD/73vvhTSUFY+lm5FkWG2YQYfk+p3BQBQVaPj68IekfjoPtmSx2mIWbHpMnW1wVnL8x
k4fVwbk4Jc7IgrG+WqKTaRlQf7zB2QLBEuzyEraalm0gKaiqIAZ6TdK3+Vk7fzrTDlePMApCw4dd
2CvIYCFF9oM1Hr1HyqfgYucFLMt7j4UrCdN8cIzubfPXDddr9z0FMDQB3fMEB1GnSQ9ScRsgAe8q
iSIw02sar4X4Pq4gsIvnNFeMWGhYW7XjN/2UZrvbdwUzGWQ4+cakJ/NsX1vn+0fmD5/yx12qhMJS
Q1q0RAFLzEDQNz5xqYyNCyhS6Lft5Jnb2KmZWRSYGiqljxD5hw52BI4laYIKUbe+u26sgIQVm9Jo
QSB6xOU4uktEkazbJ235gEtaG+QGhuumokqVT7DztBGtfADMveOr+czPXpYZCUolFwBGYsqH5Zab
qr0cYrLe/N3Wqmb6A3QRciDU1Jl+nda4C0nm2fPax75J/7hT2be4BXCjaT+rGRfW5hlFhYR+m6aN
BtSGPrA/FCghhjZF4iGIVjuEKERo8NNOypHQyJ9JxE107D13G1fuXP1zdDpkgN2M8Hco7YQJbi7k
vdjLMP7cfnWLnT5nsVcefFJiC0jiRGJciH2Q2JwNhbQdZUsbM6rSF9HTb/SCklqrDgb3mbrSJWnK
ZJ9G1pqxtn+h9I41pY/i29XfS97RqgheLQk9ErHWomxpB8KemZk+oA13EpH6CVKipDslfW1s3m8k
kLCB8gWdqbeap+wK+MrWWZGAUozyzoUR4zGWrzNbd9ektEWy6wQuTwo+VQwvSXz0ZlY9xSKqWVHb
wKBg+ojw/UUI4EsOgICl48+vsNgwTNuNYwFDz7LfbjZ1wIvQIXnMJf2eOngceRHPdNwfMs+V54wt
rPVZbe4rIINr6ekBJ7PNZ/tSDv44teGY+yuRRZL9AQNt9YZkHNGBxLgVK5UVT+6YnLX2cRI4geyq
gcIhMItZGsNMHcUJ1FpQv6rLsPHoHFEkL5fw6Ze9DDNat3UoQV2rf3mgD00W378bgpdEI9m4SZnP
VdGua+qkuP9vI2DvqB/+inuuiy1AKw85DxhLmlhODBttb8oOLccmD5ybQ4AcrWAXvr2aHEHPoGo+
A7IgUY4RLoKQgY2DaBhjCtcwSWYcIunlyLGGvX7u7ghqxdo+OTp53nL917fu9PNuvsRXaWXNFra9
z5Z42LtblOTzHntg1hqXrdRTrom0EG5Snh/LtfJhwyI3kkWsvds2uKCiYOyvbLhHw7k9U9A2HqFG
+hdS8CW+CDhCboLNfdMns7cSr/7mezj9BEH3Go0UvuT9zn1sRBjx860zJesOS/j9JT25WloQQUNd
hn+s7LvqkrKRb95YpeDvThlswMtNiAf6vv9aHIikck8lch6xV5Z8IgVkce9mJuE/0BYQP5iq2r3w
czvBbVv3Z+nscCrdrXm3lbHkrrG+zKb35MBicFN2KI/8vr0q+dtfeZYIwla/xHnsZ3IqUfjvzVkg
4K+m+3lqMjf6GWmltM1wEKyPCumyzLTH7+Ovr/PR0C6mZ2qUo6GWDDpHuusQjEd02LnKJEIwLZG5
xJGsk1sbMpK8DCPXc7gAMA6EgmFKnP2GwUDUaJzR9tWJT+P0TIZNO6pKF3QeuKZYGMpxERwWKwoM
3QCbX9ci40sO4edOn6raQn6LNMYvUvxGH4LXHFRFTRinESsv3KJfyNt03AT5TEKFMu1H0PvAQ6R1
T6MRrdIrAk5YuhX9SCAQILEMzv6lmUyeH0q5frBuiVJjYjBDRPcoiqbpMndmoHlzqrr0dF17KFyp
14QKBi4Q/9j5Ht98w5pUTOXGFi8mR3gIOYP4qB0g94A1TyPAA7Y1LgxVijjOrUJC33/A8NTSsYsp
+dsr3UHZmuWxEZ2AhKy84motZzoiVihjtBkvBJBANWAhXxDgHmC3Hi1gulRpijTKWHC46MpJYfEl
EtjgcC3c5u5Uy34YV1sZjAUcW2pa7zITRNpwZHwB8gd0DWJpHq3rKIN7XX4zXoumFI2uSVkbWlNl
0j6sxFR3/i+WfSeZu/RnEeK5O1JTMk4FwSiSh7Ljk840H2J5Pu9oRCIjxq3ekE9XjZ00kEe3pEIY
o6EY5pok+M7WCPuTkBvT/2/cJQdI1lzQaxwopNLyZHZoA4qfIYiAtbcIKVimjDaFqqvSzitqJdfe
HrOK+EJEGwYZ+CVHUcRX9ucCiYsAqfF2X1Uuz9gKVbzJFl/5xWq+nsWcUbxSm7Hr8lHs2962FHN1
rH87ZuxHomXvBIRpmaeUvYY8tWtwhY3YoqytM068j7TnoEu7yV63M2VONdCT62QqO05rffubP4fx
jjjKpB9GDJlgj6D/XN8hhAN/2JWgeQMJPAwtLIbuUQ+Yz1zbvu7G6ygSc4ig8skrNn6nfPMcxzBN
WWtclB44aefzddo8KZr0gIRYnLP23jScGfUPGDxKvpeD8dYGZhkZOdizGWT3GZKuNlT5h+lVoGHs
wRf5BZqwkPl8lTEchnf8/wwjk8CWvU+PqCmPWGdTmclBeTykWLycpV0M3VGNvOQVAK7W6ht7bIpw
z/3m5Ru44CIl4/xzLw2JU9QNJ7tNskNhw7NZhiQVcvPkrxy2OAZh/6KIJ2j5pU7Gd9I6hr/P/XFw
ptpkSayTWVGgEkGjwqdjbPOGBOzTvHUETLoQQU7vH5C3INTTPVpxgZyvzVcltGIAjGg+gbNDQc/A
8LGl5VBg1v2P8APuTmm5tFyf7L0isUOFgkAT9X1IORvFWzYdsSWl3WBUlLtw7dL7E6Qm6O3iQkpo
JdS78EIFglqUPrOkJqqZdPBwIM9o4EN7oNm63CPtSdXeoKM9EK8PmkvHA55aMv4CseGiiSoXjJfy
Ky4SowMNWtfKXuo3s0fbx777IqXgoesK6JHXuE0QiRz5t5nvw9d+pHGWEWdTNIEUSLojFv22UAY5
c2+SM81vLmduront97zeGJ8ZWpMnqWINv9HEu0m/4xIpYGP35el+E4vI+LfMHCH/8mYDYo7yl/wg
kMw1gShRhJkSVVYZri0vGDRA0G95xqZSYNFGMHQWCW7qA+LzSw3OYNeptUaDvQ4KKLsBCP5lBpu4
8fZUGK4crzwPO8Iwfkmtd4+qAuQqqbybUdt5uRavstfTyR0Mh0yz7frmaXWW9KWv7epF/K0XrNRc
MOmxepbD4MDScHDCDdKB2Ch2D0zHWs5y89R4L5RPbf7gF2CxE4eIGl7pZLSeW824OEZ4m8PTURTk
FIcYu6P5dmsI00LI+7j9hTbNjz17dRpbv5FDuE7GLNi7Kn3Y5TC2qTXEo6S11Pwccdg5TaEECn6M
sGb+B8gXKy+LeTKzPmSr5umbf/BVpR0M5LkOUWBB3jpr5SPNV/dUIS2cSnY85AQvphAxRCC98zqR
S3oCtN2L2/tWWvS/MrF/Elv/z8vIaiovcvDuIXRFxpwCxw6q3r+BPVr2WHyFP4ZUIaM3+8yiFa3s
OrrW/4vJ8alJniuIFsmv5nQa8yG4iJYT8UZeBXlZRWbz/1ovVBlrXrZzJcrZF/m5vWFusD80ybKb
OYQ1WfQqFQIPsUzK5Q+qaGWHWjUXmfxzwCs+630Jds94NZBHzAB/B/rl4P7QtJZWLJ9GT/q3BXnJ
/lsRewZpHYS/LRquGMGoxx+w9AcAc5l2mY/QGQWSbgg0OdBxEHxbzSWpSZuaIEvhyeR9trFaue59
ienZaOMZYcdadvWczwTvS2k+cJY/tDKZ9j6pMemEAd0tIwPsPHMlvg1pOKqy7s/Bc3zJE43hJnSZ
ynls7lq0h0ITao4sSWOUAsrOxpcWPSysL4eB0Sl0rlF1h0882Xuf6pTen9ItZNX7ullz55bIEbDS
RHFB9qzYP87sVwdvlQu1/5xM9LgvUrlXMMGswnvivibH5WgTbGjc4qM9tXPv8voOtRGi+1P0mm+n
AvflmFSw7z5QXJd1Wu3pcMwUe3w9ETszi+DwoZEVWEd1kqUgtYN270LfJgIY27LzeYosXx4qCUTQ
WpBeFtDtziGDgNweKQgS7vxvJvDllhQ7jb37avnovmZTUe65YNfswb2I6FbLOLT5ePvjJ3kfXXoa
8TwLKE5+U9nHE1C5Za7tA6YyNUYQB7u1cx5eBCNQpvGNEJEyD3QdeuIKs99JyD4Z01LAe9RhmLeh
wETYVqyp65ZokpCyGbH4YSrUMRflrInBtFnUX7h/nq0fFhxubjtRif4aq5SJBkKKdYraUwrM3unu
Uv+dOkzXgqYIHz/kwxMD6XUoKwFMbsLhoQaogISw66CvnejxQupPDZE1cAU6kXVl+MOB6CRdJefk
3awI0yjxOaZagkZemCRlccnH+UAR1MKPvXVSZj6zOgWIRxdAoYri9lIf3fHvvSIcg+yz8/7mfgVh
UjYJB/QteCmkzikBSSRCEvIUdzXlM4N1aq+lmyjfz1NNXzvDw1uaHv/cKq/u6bxnok0CaLwYf9Eb
X/EZPaaULcYxZIT7ZMZKElbb3bYV4e6dL/GY1towoB+Z4vbTruJFLMqE63vRaC8k/san7jk0lZFB
btBK8voG4W3sAoIvW2GGydCV6OD7tn89Ggb6+mt6tF59Z5I6TvFDBhdweCR5/q2uk510mFKiyQE3
PISldP6/hMz1iyQIHu+NzzoCGHnZSpvVWWUZHgUdOXHcxA1HeEaYy7W3cR2qGgc44x45j91GRT8X
GVhZkUL8rB/S/fVNrmA8GOSVe+R/SWJ/tUJmwoL/40HlFfXiaZm7hjm3qNSVNyGb3hadFPOHwqWl
BFNb6L5TeeG9n5nbbHJBOCAi9c+5MPu2BcvpGMPxqfGZ3c6HC9cDWi+0mg0jCj97oHHuALMqI9lv
Lt4nxKc0LYWO+8o9nPj7H7IfgkJl+Uf7730y9cE3+HLIZqIq5BIEBziqeWs5OxZPVi6hOM2KybMp
orXxAZONhdfvxmkQZg5nnbv0lq7JJ+wEpi+g7R7H7nBOkmK+38FXNk7ZBZExpk4+97jEnrnIx4ki
q+JDwSdtEGLWpw6VTFqhOZbtRAJprR7vH9HMLJTTr0Afwme1AwUa8lP9WBZvmfpcJDhdnuQj3wbh
COCLksTXDfM4jDdzSRCwCeVhRx2MIIvjZmEE3g1crHqEt7EWYc8gPnTNo8Z1gq+ejJJn26mDw/r2
1TwTmLpBVlepG1b3QtZTJ/yEcVbBDNjVJCdv+RrWWecDxrhrJTALYbVBcwe3uOMr/tbFZ1Ay0cWP
mGIcT+6nxFjDJXStM7fQD5NgJlo0191RZS06aNwxpeC6IkAFW38bg1QmRIrU1/2T/KI7k5h0tAp9
UAdyx8UPEwEuEOKKfm0ZNN6PlciUbrXYga2x3rcpzycR81R1Flv7j+OEHcJuHkWUcoHR87jJ/pNT
Xu6kqSkMSoWeQpdpYKdck0FI25Fa9s5is+H5fGGB2Vaf1yVQsQT459xz44y2Kc774h092tkMcTUm
WDjnrx2yCiydNvqfZuNVt4+xRhUkHavjGjOaqj280+w6q1wY2TRhv8n/c2JIZnW9xBxFoax73Em7
9Af4OKmH2MKztCgkn5MKm9yMhe1Aic5XwJEAVDNf+reRBz/dFlwxOVNYl1EBdoUrBxFhZZQBN8rm
1RGjijSKn+7MQTfRGdWWKJxm8h6xGTuYmRRD1VM+ms7pHwOHe8f+EpNwzUIJQoYKICxl31SJw86U
6hgcdQ76mZiIkf1dS+pKS9wrGDLlyZbA//X1Es74i+M/gdXQWa4uvOGaMFKper97EB9VhJTzxftV
V0L/AWWztkjuOrBhfkRu1SWG//R8zFmeZqoe5B6a0KCymMYqnSyUK4q5gxtcQZHrKNC9o5/gpNSU
FhPxKjrTihgvG48LjY3W/Cwu2QYOmeH3TjlHdNiZ0KyLNWHK4bw81TAwgFBx9jAfkiK9QKKv4FjJ
uJayDw7CILkLAt83QD2TBlXHp1bglY39NycMjkmcMUk7vergwGyKVrP4wRdpY2ScGqVegZwOKwH5
Vb7GbSpTgSDcLavYMJdx7FKXPcqYlWRkEGBXtTBO+TH2WMF1+4L2f42Vpi9B7OEEOa+mhn7X0hOp
PpzhcBfWpIo3glMs7iuyjdBiN98jTNaGjGG2T4o2Tue776c37Qxbo7bU7CnbqOq8+vKarVNiGHCl
/33t2Zgf5H/EUIkDGkfC+h7Lcf818CGkFKiOQL50SYjsx/IQkYRQHhnV5Lt7nO7xCQDNNzaJedpS
ltPuWg82iLjbv8aDRDeQI2kVXI59h1CmeloANiBbUDOiMku0bPHA07SLqUghmun6bY7ClXalTCIx
5d7s79MlSe5HH7EvElCbJEe74sZtb8nf3KqAjXekWguPru/9P6GXZd4hE5o5AYjEbcMdTjOnA9Jg
ehqzDaPHqk/zKM+FExaraq7LK0rBsor+HwiwYgpL1mRgA+lLQnP4pWMqqrMzijUsKa5uNVe1kExF
FsdkQca5LcoZy67Ru5ut8GjRayT2dp9wj4w6kRtGZuTKEf7JSUfZiTbCH/QLYEjuD58ZJQSP1jd4
y/Xu1njpSGgDy/c9TF1xUSGKJiBDoFLxWnJhR50ru5hRroGpbO2frSBCvJ9ZiJ8MiOduT2lGXpgW
rkEqzVlGzBl+S3KFGxaiqsu3rteGHmvHMsplC+xck7LFFbp/s+cWOzLzAUrn6rc0NvAsDSbBxhxc
aYsfKA+Hk2E3q4UorTnTbXLsYaJmwzllc1LfiZbVVd6xUva7i0yW5k+TDT7m0+8Eye6AYNhz3M7X
C9UEUQAdN4iYxL68FmiApvlQTPfhJ0x+8jTjvYQ7IruXdp5lL3vB1iQvxIWMRFY2VYuEHHWqj0VL
JEnNPSu0Op10haWuVmlgzPqatNwEA/01+BF81bW5hOs/OhaquujWxHdBsMbFz9sZUXbzG8clfsun
XL8rmmY68C53L+nLPWXoqPs+rfmvQzBDYu0XhD2OfbsM4f1zPGxHsQtzZvF+zYiVfrQdxm+/18fb
ggX67H/0w+krTiJBu+QA4Z1df/BLVmmmensBqYVGVb2vvlcln5Y4RKmRrHncHTW1IjgmrLdGhsdw
41+tt8p6IM4xJWEvl5j1Uu7eB/SY8YmY9/N9/f5+3yjA43kJRKPSl+/xieWbV9Sp1MWGmtzD8ljw
gdeKDeNQnUqBAuel7XuyO7w2Cl0Dq06DRp4o1umWNNPSb4Z2USegG+gSyVgoIiG24u0PR2npzOxo
2phbgW9RBt8pzMqmJ3eeyzC0LK7wynIvRykvZgXlH4EmDyn96dgcsYa2e5sKmywgfVR8lbXAmeII
04aLuKZADdjpRL4jsbohrPpztTv0x5Qd1ZncOnT29Tnp74YCvnfwNUkCg+gbJGSXSF/onEina+jN
h8bh1qXBtIxNo8crd9516VShfPZ5YbCdsdNhPOxlsd+z/jzl+aTWKw8xXJZzTBNb2QxEJjU7UR4z
oihEq5uatdoQ1eYJKqUGZmqz91epkTyY8u5nPEIOWup2nJnhsI3bsFhh2+z3cYWfa1VuMoPNiS41
V+wTe6tq0elyzylAUQR9hfHWpPvZD3KfK0h7ZroUS0rhd9mE9NbUJahAxPP+cenUQwK0axtPOTBD
12MWffxMltimGux4rvCHE+QccLPzvGaha4s564kVuY3SbbS24GXy/rDtk8OC0u4qC5bw4WKqieg8
6OgUB7NUtf314bgwyAezTxaERoe40tOWyn2wNnwPe9wsXiAZXyasbbjuooAYB8ea6tsNwQiSFxnA
m6OzqtzuJmC/8orAjJ/o2or1gKtp5P85tzMbaTKhE/1jP0xgMbx0OXGfOdUWqTsyMhPqwfA2kudI
xIm+zj9l6kVXcgoYkydzJqHAzd77hlaPgcL5a3BWNs51SmbsExMHTUnY/ixm0nK7MK8teQx1p1tE
f6aDHX2OiiY2yro+I5oMzOSX3LBGPNCVNn+Eb3OJcwJLWdXW1cQIaXFswXrircxCGNYSc/cEf59f
IEohNm0LhGLapOb3pqZukv5+52vdhI9qP1++WFgu251cE4Dyyz4FUJIBmLaNIa8r4IX+qeZb5jaY
WbaNrKMQeEIesErk1isG5Ap0uAJmkl5T5MK/bJ+LkeVREcnWMRqIOkVK3q0+Z2Ex6r1zlOLDPXxn
mPdgUutdpcHPxMnO5+kw0mTDjUNZ/M0dpsxe/GM/RnTRuhtAV31yug0BmDnzAL8ngylzCskXm7AM
/gPVA4JdgqsQyWwWn+W72WWkShpoC90Uo9y+5bw3Q4ReMNsJXQ7v8Sd4rV9JoopZvKuX95Cs6xzg
hbe28b4e//hgO+ypUnyEuBot1rsgv0MUBoVl29lsBr1xOePLBkpqkisk+wG1Q0SK4QSyRYTYdgbE
SRd+yQ5TmXZWtu1F+idTykP1w83F1h4y7m122BnYMXGPEOffKJg17nanmJUs6+thKB0zzqOULtBH
wuBLsOS9BN6GpB02MN8mvIpzXIbfT9NAu7kg28+gmMkXP2FaGX/x0swhBohSrKYLQyOt4IrhtDLZ
WsE2vH4H+sX4YEwyMB0JJngKrbgTglBdzOmFj+TCAams/J+tRBsCQmNI+iNAO/xEMzedR+2EyGPE
5F58Q4lM34n68pyXPzbrKppWFBu5pgM2F3hT7psg8ZI8EISoyUAjlHiibks7FTOZYOFMh8NyNkWz
E0/kMgcKAXHdASC90umK1VHO+08G+JLdTisecpDBtqPVkRS9sXxM4fmJCjDylZ0i9XKbV/E0rP3H
UrGozAdxIGn0P6Q4isyhtUKbr2msppbsyO+rX4tpPWQT12bw/plEYQ2MFURmO1HkB5t8EWD/rVPZ
OsI9HGfjm2ndY/3TzJ9AfSJfPYg6T3JCRuMduzVXHaqOpvJ3AqoQF9bUVq61eZLM/UuWqVSLkfVK
+u8sfvCXG8CkO+Ibm9SnOqrSpfm5r3oYiZq5EVT2eMuWJlAjNWDnV34m+/j2sE5lUKLfgh2fDQp2
fySp7xUHiTzQRzYTPj+x7GRkfMnKFk8W8JodnwKqqoHRw09oG3rYujiArJ96y4cUDmg64y9H8ALG
RXWiETmsRPhaiIeNhsFw8etSFvhemB7KLZPev2ZChbbA6LbtLOQ3NS4Tmiw7tE9CvQvBZCHVGzWT
fN0X8KSN8v6hIL/fv0JgyCmK3uHurGtxUdbMJMVyd/mpWTJa9S116dMGhwa/ZwAUUuXZx44D2d63
LGqf5j4Y0Jt6dsf1uVl+rYlOzaklEFdlqGIR//E1lONyf7xW50gwhmDNhMmIaBr/MCQu4q4FHf5w
EfOs8JZ+W5m1zq/PnYxWOFXruyeRtWw6smels+URFsVQSC92FjLIoZgzy5zdeB3JTMuxxPr7VCVj
4f+CVjuui1AmuBGVPFIsi/mCHTnr6ssnp/4d9B+XwmjS4MbXjv2PuJx9Dq2KYibNMpo9AsWtcKUC
WUkyLJsRC95zEbDmUgj0UGPtUP1VH27OOlazyVwquboUmHz1rEdy87LQkUgl/sZaOrSr7U4GZUqs
RVZJM0/TkxyJhj+unSHHW+cxb9W4Y2mGCQU2tXNnxINTQ2vMUQJNrwZ05KXNteIYgKGP2A7hsLBY
5V+5a9diXJJRHVHscbXy1IC02TsFdR+Y62u3PAp6xueUu20tWWGDkt6w2O8by3YPhHXc5cOkhl98
QwZDpuq8zDGTznze/K9CY6794EIxZNJp/GDAjGlOve5wLwtRzZwp1C5QgFmD4JkHpSx3clZuBeDu
4VCsexiENJzpAgaeBlZ68V0ueWtPBaeaW5uN7mbrRafmoQA1BNgldXcbHoNQiYVwQEcKFw1VjxS5
D2c+CT7WYAqF9ZNQ5VxyrtqQ5uHVK0UrhvJSCD6UfANyW4Rq5utIOXfXb07Iq/pXQNPyn1f6Hr6a
zi+uEg/DD+vhq8KwgTWapbtfcm6Jn9gycvPa/YHQ1avn4CEIvhLsOmgrUvt3lhUBCG6fXGyS28uQ
ZevUWoo9DlXS7ZYylzy2PoijncmqnUuadGvE1rp9c+UL2x/HHxc3w2joFVRS45oJ6VXgbhH6TnQQ
isOPipVN8tjWkKSa+GXblsFnvE0uScDJSN/w1s7CY/AZowYVZb7WcAjhLsS97Lu1L98R4fXneWed
P9aZgcX6bjQQNS8hhHLF3/aWB58r6Xsyit+5lw01Gywvz6Guj/9MOw24h2M6KOcwktA0nhOFur4H
eCAH29px5PVw1GqX/PQBohAQOMvn+AY6g3Kp7KGtSC66amMWKyDxHG7ls9hLu7N4a2/vskqvA9KG
yxQECn6Cn+4Y39VpXMMtUofvtmCq3vGKA8ZAiPCiIX3NEs/5WrCR2XSdz7llKO4C2xKqtRogYlg2
YThA7JvRwF+39sj1FUjr8ZPHFTkIAOKJWs5c9lftvmZhdQUHyyKaGtiYYKFnDgRAC9Dr7LRNIe7F
xQvZpEMR0wI75xsIAGqa9xzyIoiZWgIHnVTEnuf9BMRtdt0XMli1e7J++rFEeElSmUTx5ja9O54K
Pdh2+kFiJShWwJAHy5ti1Y4vuRNWHuAOzeJKB5OYK5Nz1ymiNBBOqerLLVjqapOszeCyVo5FMPy2
TQ/x9lYcT4d8r3aG85erHVkNy/gZZykrucz2kawpCFPVYa0ZAAtKs2nlXUnKplrvy3z0TqR2G/uP
qLGErxevrqFJCz+2bOgUEh/4WdzKxgn6u6Kodd8g2pLX+QhVR9eUWxwa7MpB4KUPkxdJ1SbSRewR
b8DkYq79bd9ehu8mvdY5FbyzJCHR/QkJ+gfVKgqSPdDGPbSovr3D4eCzmEVlVpRKZOMrmZ2NBHaG
C6iUSKdpxXry9gAxPSioqWr1df0hH/2LaKBrgNqQo6bOfvSJYH25ZX8RYKAizjuYiIjWR6TX5fHX
IzFpnukASUy8Y4jI5/Dcl7gGjLgz7c46ErqTw++p1E9sbaC9yQRKdaGMoM2JQLZZPyoogKAE/G1j
cFL8IN7+M3DnO+VqskPNhaXPEDQy1qKt8kkQem6sIlsCDPdJfp8bOThmGgfGOmm0+f9RxJy3Lum5
17EXNiJ1Pl3y7FeTAXVw4PbWO5NnP3SRa9GAwGmTgkDB3voArMKO4f4Kc3Bo6Z62q1ZXt6QsXYVY
QaYKhepa4Mh7byAyy7c9IixgBDP2xBBuWW0oSot0gHW5kJdhYgBF5wkhcA0ICFpC+ghB50d68dlF
5FAkCrVHu+3HFiBIGGGF2fMCOMvk3434FuyJ4N5tk9xwMmRyrNYANnfuYJZkkKUHPMxRTYEjBsZq
6XoL1UdPdHDYx0PmlG1j13yuLlbfgpoLSmL+yo+3TJN0r+csvsRkhI28Z5nw3bqwbnaxGv/O89mH
j/GBzz+QTGfI/qhtmDXye3R+Hi1w7hHEmg9J+ns28iegZ7JZfOJ6RZPyYwaP89c6k5M5zrblAVwA
LbKh0zyS9GoqaS3/wp4PMsmqAhWfnI1pzeZMljanYiZgutG7lSaqqn8eHy9Rl/q9/1NKHIx4i0El
HMvak2snPtPH9gm/jB+3F17R9c0ObXURehqpnL1mZy1lmw4+1StREQMaiXWVlQQ9fMuIcXtTwHVo
3zRS85AQckaiyJvGDyg0cAShz6zHCF9BtdqlAOnFgCCSciN9DRaS/uTgcsmM9Q/hGRe7hYA9CUT5
TJygomjrkSYBPY2iHpdOL4WyYt9ru/bnolYhdjXkO0YjR6Cqqy3lVwe58x/mI3NtFng7nyKJjDEf
fRZoCfGIm/Ynyw8drA6S6zmn/A5gtkGrxKQz+FQE3uhLeFiZUaJHp8Q5gJspzUODp8iqJx1hQk2U
0U4y9RhbWPyOtIPzyHJ9+j/H5GHho2K5E0XjJn1wmb70Maei9Uii4GFF477xc9lK2d8GI/OtG/Gk
FR1QBOy1/XeDFsehTK9fDh+H6ET/rT/YDVmErQsoPcn5f5tfp6hsnvjpKcV7YSOm96fHWkj6mC2h
0MatGtf3DeAYMB+iMmhanaVDGGfWxMdxO/9GQ9m7Ax0tnGtmEGZyGon8b2CR1n3r3nPPeN+5hpAl
682c2o6nknmmVgdPzfXAlOoGWSNJkgGO84cSp1s1Np93Jgat0lRnEfcVchD50bQwGbZMD7XcPbYc
DDziHUq5y8jJXgj1P7Jndhrkn4hjhnjaaTkXGTtnSU/1f7wg8lWy1FPf1PodYVasacLiYMvUJdbQ
TcmJSpbc5w4PHq+XLZUHFFupbkomy+BoRavrg4ALgbrQbZA3VEXZeRcXDHsSTz6mkCQDhysFwb3F
5mrhYPRUss7e4LOAY24Ph0eS8SlyuccaiH6mraU/RLOgACr7z6gQNUSxbVr4laZ06BOI4UEmd5P6
+sDaRPK2/RscO5S5XOaiRptbLuDPTHxOgBs+JjxW46U/mWPvbjZnlScvjZ97qvnS/fokJ1lM0XkX
crLfQWpHc6P0XOPHz2jyA2+Dudt677A6JUro0JAwSNDgjc7sgNk47G6JsWHQhT3x+w6ZHbSFQ2BI
7nSPuOIiSPEDsKUgsgd+tslpxmxu1TqnUPOsT7DG1LkmAs0lpvruo51p+G4JaEZITnpKDXQUlxAn
QnQppaTSoPz5BRGR56pxYi1GNOM5JncKBYRB9XoAS7LbOFuGjZ/AbOPUplmPK2LoPlYCCDpdzhdk
jnmWoIafb1UDDxIWsrbpsRtld4/qS1wcyAEg7A+YtyEy947ygsrXf+ZSynRKu3IoGf5v5V6KpUmr
XnjI6svadLawtKUyTnBw9O1LXRomR2R5YxIYWwsaDfa+0tFPWB9FpvQ7vCYr7iPqlGgkNUNpyq3W
4TsJOzmGG+759zX0mVBAzM74sOCgEtwZoG+ANYuvYA4eKAu8QIaV8KkyQYudOkv7TC1kSICy9ZkF
HZZ5bWcYnoo1TPDvETYH/Neq4ED1FAE4ksTHOpoCV+YacU8DVeiCk4HcsQPv9ZaaSxmEZITngjzW
b6lrefVOt0+l9kZXOAwrb1LaO6GXMfFYqt9mSG5fKdVHo80/E1w5aP4/X+nZD3p2Z8bJ3BAzijko
sdgBeAgk6RAdhgAtB9SSpFOA0SRt6RgpJ2tV0AEpajg0G+j9YJ9PbjZPNV3QQ0q0Vwy10z4NTD8c
t9CUhTZnOSI6A9bGBfHRdNf4XcJZEdV8qdrpQRhwDJP8brGLePXLU7RDhVju++5nExF7Zj8Lbe+2
Gs0+2HMZ3xAIHhCMod+WttlaR2ecAVsS/eszf8HVxrvWSEsLqz3jJwssOHulYgJ5f7/qpCiqCThI
D49/tJo0LGVZn38zN3RbvnFXNXzfsBvRIOu/Zni3bE/N954xFukJw2xyL3nVlFxyOR54K2iIxebw
G5XOqu4/I1LBXIA5OibE01irLuNfth9zegrrGL2GjcFh63WnMqF/wSeYbw6kXjdUqPgq1a9J4vLD
K6ZlxKGWVJGNRAuDx2cVC1fs4oX5AqF9GWGx1Xa2224bmj9yYzqN2aE8wV4k3MNIzjbpTEmBY4y4
ozAKzYEgThT5uRRbxfcPkcGY9K1c+kzRwPMN82PCWW7VepkpsM3jzDAMS0JTZGch5rkgoUUnWjk+
3pIvrWjtz/zCEzn2nQd+LR9XK2YEuQLI9bkECiPBAeuI0wXs608lNiiMWlg1GxyaNYZJtIoK3Mo4
+Grbwgw64kXFz6JMMGnwUd2YP7EW9QTmiBKD+3LptkuvJdlIVhkg6O0EPBvhPU5+dYMCfaa9zsFX
QZHnNTuDl18AafVrHWF6rBllRIOpEivot66exRlL5cf1mntJrUqQqX0PfmFzT2xZPgd3nPje+iIu
T3rUj5Aqt6cv9c/J8IuJNOqFT9FJPF6QJC1Ej8hbiFJr9we7scxK6J1DXsRb1/PNVGBeF0z5yGxI
Zt8zhaStGPfs+mtSGC4AicSY4ROF6V43GYGRheA70xh7wcFVx7OjIHnbSU8e0Gk8dqj4rkwpz7h9
VtsOXTOJQfwWobdA7Jx10l6LNoyRyIyiqlXlRFMYGNXu7ff+KdYohVQsBRA8115nTbOWf/fojAjc
ikpT8UWVNiz1co2E9WXRfDBKrw8WW8QMeF7UD4WkzB5PRIeqoy57Uz9X6ymQEDY243QhJnMMoII1
t7kJWOvt+76zNELq82LnuaTDO+3QBp7iEAGQtWgwDN7kBbx5EGreh7dYDC4KdJDP+HgmHdeHMMqd
Zy51eLw6UR/rISY7bjkm5FxSFG6jk1KM8M4lvhze3M3JUfCRgdoockNRn89+e70uRv2yicJyur9K
uUaRW4fohrwflxmKF83fnz5+vALAQ+3K5aTDD1kcP6vxTVRw2THNujUwLxvVOLU7o38AxoLYjyPI
kLSQTTpdZTCwT4WbjtxlSy/9ieJcm2OwM9u2v7bDRCHxcWA2yif1bVPO/VVo8Rz1YWGlnQzeKJ8E
W0pDir9YTu2edKnl5rEKSG8Wls7Yqz3FYMHWBDe0WeSw7H6KjsHZzO3SOw9aHloL0J/t9z4087Xh
wCPo7sj+8ii1C8cYvn1eZg+xDQoOid0/hdOtiUrZa4J0xm5mbPtvqhTRiI8NRvDkYJwLhZ7fdTaD
q8cxRSXhgqzz1C3R6s/kJEq04Zp8qqSHsZNdiciVpnWTN29MnTZv/Cpz7t7klj+HFFKmS4ivjXkQ
knCdgz2kJ5O8Izb4jTVzBJBhO/c5sb6v7uQKOwuqRuMDtRz6B6+kY9K9I1Vs60MKNL8deqcW1l03
aHvOHXejncm3Qjq1BtZfcU6zOe4qYKPL4BWrStqMB53uV8tc1Jzea1XbPKM9Ip79bKFBqACm30uh
eMC6WyCvNx/WiTUXrswLxmTOX8GxnxIHysz1NcQMveSE26Psfawr58qe+O1aNnefcDEJ1+jaPMb4
4ltG1zsynXxcktGr3mbF9gA+wqMYmUSUqQ56c072p7znosd8JUWDhN/LQYjnPpmCJ+UjUMuSEMpu
Vk7XegOpJvMBmGscbX+wGx7MhASEtPaWiI3x9Nm620/pQq3U1M/KAkPOUBwBGV1wBvE3xfui95wr
xt38I2YO7mKl1bP2Lh1ttv7pOBqGBDHKO5d0E4r1HoK1VsW/gorXjSQMFEos+vbxcnQnQTV/i25o
PsthvRnQPTrwd5Q9qYA/c6JB0SRegOyHT5UWso6ce4RK1tGrPAHWtxPnZy5YREzQ45gv2N4/QS4i
qSKlx/12tW1GGOoEtfC+xSAxX6SNMDRAbPXFoyh410mf0IbfrB9fD7cOk5mQJdIKOXoUjLT0e1qU
3J5lie2qftzCnach31gSF5mBVd7C/kWgIGH/3csxRRdABg51TYm92MMhn0tb89PEFur5ZOo5Mi1T
ymwzkcLpOAZrUIbAroEPeJa5lKz8uORti1lm+KKpuX4zT1fx6LSWTBcVmreMo8p0WyvjNNxlLQjw
B42SaONW/SUK30r8kk5Y5jx+ZYkXe3U1XwFf324+9c1umu1Ku5m+Myb9ty7Wt87Pf632qOPvjYoN
qYM10FEAPPoQEbah9Q6oKAv4GNHVZPjNrq+moMGgg2suv5DwdbvhBtei2XShZa2A2Aw221WhWhVP
kyKbokXt7rh4C5HBDA0JuW+aJUCoaM80sKyYDd6dTYv1iYk9wq5JQtMgycKuRc2gMJbEoXXtXTGz
sYxOsK7WkBpEkObNoTFlwOS6JcArcAqgpW6ckkFiajDzeY10KNi4kDc9KUND13HuTfbyi7/Ft6I2
BFyZRT5Cix1RqMsLdET+BFkfBfv2lhQoYurEsw2BfgXF7jeRshGFh4JpVssp7HjY7f0+JCVGNuSK
P9We29W+/S3A7ewuQ3GA0Zw3kJSwhtjHiCYLVAnKDYlVsO//rz2lEDBDPKDMJGemiGdyXZBkiHbr
RCsyPQiyOgGHYru82ZK7tk/h0aqPuXEGkXlUb3d9ucbmy7HiYrvJWUqknVdB/pJ+VoVAPat4u2QU
CIsg6yrK3X34MPEVfhP6NlZez/r9N2hohNs6dqm4hy1b3kT7MGppgoqTnopDw9cJrHvjdQff1LTz
NuMWyPdI6DDBd5lYhA0l38bK5JVgsGtrpnlPwC8Xb5IkzHw2WtFzr4EeTVrCTtvE7LVP6tMoIrQI
E7FB1EgaPgVe1f0esFGeW1CLgyltYZ3MeIClxkcYSBCcYKK1kzq6sKFaiZu94/aaAm1DndhA1S7p
11yI0+vv7GiNNCiM3vIVkExC6RWAifr+gkA/PGl4oq3cd+SPHfnYfnOvNWs3MQ093Ff138mauPER
bjn2OGdQsn5iEMZud7Zpy6O33qmzvBSN1n0qGn9b0p8IKQm6oWXLNWsCx4ey+AuGlYRT+DRKs8xg
/ZUmqWM9q2nGc82JNPpFUoamZp+6micS10zDLR7oFqq78ZehhwY2ypq6wnDR5YNFdsvRTOhm5Ijx
Tucs38ho/cs1FbuZHbWG1wI+UJSNO25iGdNZWSXJRsFLeco08x9JTWZ2G3GW13CNkZzspVQQu1Uk
0OBlRk+E/n6nEBILzQIuPxnpKUpYaJMF+o3tB3zNpJqmzcIPIZSI4z70uA82okn1MYUpl+XuDjeV
CN4sP8VF6d0Qmssd3fl3z0s3lSBDRqSyPwXPTVE5+TbG0Dr9gBEv/0wgfOTjNuAIV8iWA7VQpAZD
KNO9YDD3KoWM2LQWgm5bolVVKjetSq7lVIS3sGKnmdUyH16H5AEjYIwFwChztb3c9xVegEbTCtW5
UhMJvIaxgDtr4kcrA5cfHQ2Q2srljNdJJl9tQPq4/JXBvTFcwCN5Uf9Qa1/cXKKyblpp/VUKIEqX
bE8oFOAdKijt84PhOnEKcHtHPdgO1xh8wWzAVaeJO3VCKmR0ayn8oYnI7rklHORY9W8MaN4ODXhc
pGsFX7Xkn8ajh6QsIQKD2eaqIfUragUhjUimOOFueqhFw3nkV1nsYiP5vzdL5/uYaBv7flV3hoYL
Zt7qoL7kdehijjcBOHL6as92QOd7Io3PXVPAXcCjE7zsiKlRWbXqasyD9JRM8cyIywQV/4SLwhJu
SKrPgFNJNa7D4os18Y/4WO4CO9QAQwJNmgUP8ev/tkm/poo/HE4g59fuAmEbe98J9p8C/9VKrlhh
r+mnwnhcKPSs8WAqM37PaVuCjTB8VP7XASfn7Nvfl0zBSCv7i242NxgERFpm3NS+QLIWmT2X0o8w
cqooutwtJzaadZawlXiIAIMvPo0UOifGO4AgnyDTjG0jYTgLcrZvTCZYND+e7X49M0wJcjw7n7u5
S5HxAGPjC8BoO+jGtP6+swW9H6cJdD4H1/zTUfupvxBpsfs32GYHUj2XdaO7KC27rsjserEESbmH
13j7YptkaFB33lvM/ijrp59n9mk184jxmyO6KWI62XpkYP5oqy22oGzhsaTR6fmjk85dwp+AHA6R
xXoj3aROGgw857jKOZkXizDoBxwhpTkOOoObNHrrVrR9nX4nBMc8SxZf/PlJzx9gUneDcWqOjv4s
aljRM+5wWOUVOwIYasjoxz9oZlSm0Wjkv41qsyp/yZNDNQ4HXD2MslIzrTgQX4lRBfDBH5cGF9/5
fMdxcumjMl4z9g6C/PcG2+p1gL9bWCn3YvZ5pTmUAFuEKr0S6Gb/D6fh5zv6Q5IOMpwmbhTSZmzM
BYkKZT/rx7veGYZ0C10r2BCvio39hAHZln+6NltYfpcwqYgU2V22xeH8CBy+NXyIJsNk0SJqBUmu
DzgcyVcNlW4c1krswQkEFsVdmAZkywE+8hBx1vO3OpAjOa2cASr3jNeap7m/DBADS/5m5hjVlfOZ
r+Y11ipJ3vPXYf9fRGSQBLG7nbCDSeJBMCjpLZKfhY8/iEBF7r34VeRvzE3WuTfJ8PGfQ84IcriL
3BOGd8nR/iyQZYnyprSRXeBIOBZHf35CltllL+svQARA1H6li6OqVjRDP+sqbO9misqTXM9A9H9d
A1GSb7Aac7hN5uzlBw/hS68zKwJTOST9TmnjlEigQ+QBmK0WLdH8b7LxfvoaDkCZkDIwwOjZQ/x2
B0I7S22cfAXPwUH2FD/Doq1mR5hvYsaAeqq0deC8tuMsBzci7Ao3JgvuidbWf+NTltBekDtYHKGS
IRlul20F2wimVl9lnXdNkfiiRtRShlYmXLYliIPU6fB6p/lEK6IjYSnkfTzB96lhiSF6qt+aYYQ+
Z7XkbBeti/ZMlqCZI8eQdxP/QybcuA7X/2gmS26OconT98ZXk2DcTQ0Az2srXHuK/QEtxds7aLr4
HK3UXWIWegvb/KARLabDZIQcmRa/SXiuExz+dd1i2fPgNXrt4XQiT4l22Kj4JXIJ5Q5089c22uES
v02tv+xGA9RYV1JoKF5hHejxEXjlJtaZatrZczPBUQYezoEK/NKkxRp+EyYpnRB/3Kbgcj47HG6D
wm/UpUz0zsjq7S68Ajn012x1RoLW0AUldMhT+VC0eRFQ537HLXGU9FiD0gqbCBmd7Y4xU0sXZP1a
XYSSdQRpXYTBvpomtf0J+xCEOR2Nc4H6A4u1T+GdUxK3NiX27DGLs6srxTMgfPOEwx6Cpqdy+q2K
N1lF9aGP9TeRo4sLOnsmL4RfETQPtwXOaOHwz9GxW26QANuATLBqPWic+0ZgYRqrXyojaxy7JFHR
tXAOlwsk04k1AYemQZCqTNtbxexg/bxOr6zlOLwWGk5IsLEiBYzdipGw5w/sWTuRxIoQOiPkrzGU
wMqwjf7gtCNOH2hx2fvNkRu9A4xk5d/xk22aIMSOvne0fMHoYy3lesfZGeK9KBtdl7QeeyFtT1/q
K2b3xyox03iupJBQrhcrUKP/F+KvaofGe6jAo+tVM77mL0iWLSIi1yHUM8t4eMcfFcGLW5B9RYGt
bhbF6QJHMgXA84Sdw8ZezQH25ArdtAifLpv4AVHNrPBNHGL4MaULdQrEhFA1I9WchPApK0N6b06s
ZoRbqj6sFfdOFifqFqsHcJTFG91DwAK+Sa2BduCP09VarcJOCK0Xs1ZZx0uOjGVjUZHmJz/4p+K9
IKosaFi52NKHzDqgg1GYyjBoQTLVO4Pqv35DpqkayG9KOPM0v3xSyXnFIAfReo8QRo0FzXHz37KI
ZfU4Pb+1+QAm/zkqbz8Y/SQoUNmhCivCIVLAOJQgDyVDNywv/o1vHJmBbFIAMWnFjlUc8j/SGjUZ
raJCii9vH+KeTBdwz6rJrKgSHny34MM/Wzs9OljDO1VxFta5Ez8Mh8sigf05SR1sHeAGFTvOyttF
8O9Rw6wZGx3UFtxqOKhW33/tUqCduYB8NwWkiq+JHL5S7R3dhsr406lNM+nJ2/L91M/qfnxFkntG
YWLVtNWpomi343ZDhGBeXgyXQHqtih1VXAAiX5qDiEJnVIyvxSTKOav+QFKf+gakxhoF/WbQdrWz
X2j9y1dzWKeIxxO2QHxiuSCHTS2Lv1efemvvYM+4d9WUefamW+APjv9tRAc9+cDunEw8HHWVGwae
zSxSEpqGbrzKE+iUm1EI4EAArhbvZbi9dOgUNkPFLKeJTInH7aaf0kUVY0aqtTiyCb4Y4ttrRAhX
f96F6hyF1acxGB7lnwRDOYaYER+CD4eOp5YvLlK/AxIij25lh27Zw48Tzr0jtwnjSl23Msultgme
lNPUM5PgKntTZgu4s3oxbAl8L7sHxRUnm0Myog32fy7fm/rzcImFzezhQZbDnBmdxqEqBcdIQJUg
WDdZ40b2gdZEHhoIQdlQLRL/nMiKnSc/I3uCnpJmunw5qoN0LizcGuSiS6z7HHOfVK6uny+RPGEN
1eZJ3DW/2UsFx3wTUA+MlIYAXMatNVPxkAW538OhvzmNLH1JiEZ4duwJmjjpYYHzZ1urCoznv2XS
C2CoBlOwMLejuq6+51lBGGG691+LFXpwoBzBoOj6Usp9KdeyWdRlZuyFjTHyt+XLRBOWywD/WeCj
dqEDLr8kOo5wz9BdJRhj+1Yguv7yym5fVr6soip2A4tVuQuO2uD9uKf1dTRxdwFvrQ3Zt8wSDfDp
OpUvi8/pTcka9F+ip3YmwtUIwsHU1PeIeaBkyyZol9i95h9gHmXhCABMXbOZ+xIuRWhD22inZ/OD
dJxLMSIw7NTrOnXb6QHCxGRanF6/0dXRKKqeMclQoEDzLselYLdTw51D+A+QLJ29G1ZUTstbbJqm
Sa9UKfEDZKSfpEMt2OpEPKRbEKIh96aT6OsVZuA9BjSu0kzSlr32heAUTyppwOv2CSkwVfpST2GB
gduvionmiuxH3ppTivYLeLo7TZe0z61O53K77AMGM8TG4ncyfX5lPaQ3ZZ6T8bwIl8YWSbTomCi+
v+w6OB7z8x8elWhz7DTgmy+GnwvNjuK63zOETOjcZphKzjKYvVYgG31wXyLbmFNxEqCFXLB4ibb2
qX+ize3tCmz+LihJ5pv8/WoUEp5fTzHfbb/erhzX41xXWSY9MUjgwZrrIAc/IZQ6ZSqkx6pChTbc
WMxpfagMM1hk7Uh9dRylXoZrmGXjOW26DhhrLDEgz1eEg8zkKCw2mGAEe/EqAl3iq8qbtQiqNDYB
MZWzeKr48hXiPuKNqYrktZodbE8pJoPMI2Ukbwr2QXVmsmnRr7QMa4iuyHz8CdJjOHd+FOT1ndoB
FRoYUQVExeP/YehvdGmpOdCynTL50cNiiQVCUuNH3PD0BWB/r+rpqNBwv7QWsLpyKOEcgjaFVoC9
7kveXLNBuOsmZTldL4S+UcEjyR64Qwt3sNvaFYx5Xs1ovSfl1mWeAAIe1o52x9cpIAmQ7ZUmxB3z
yxsy7tx6a+4bYpiiVkg5X86cco8ghqGffyqnHfLu5VUMTBQ01SeK57rg2bzsn4glMj5tpUaZ4eu4
kP1I9MdWs1+1ZSVo0CiasqyNZ9Y37LKWx92VtZ7yhfegtD6qwWHb5kCc/jvBeIuEFyk9Uq0y4Lz0
+GGbEHtx0ufZ84T7hGfw5kN3U7tuRAm5v+a3ic6aCVRE9cpzmcfSSEc/klLAI92muNm2kyU+DEGc
xtcwBzov98Qv43cr7jPR4EQFxj8ycHtMDY4f3+JoFns3qB94vSIvMt1affj6siXjn4e7A7qdU76A
yUu3n45wlh5TH54iM8JAoVPt6NcJi0nCYcuZaDAOFa87j5RhlPFjZNq6oAxHZCJ3d7gnYiHSGy50
yD5XyMRzcNjgh719yjfh6N3zylfqIWFKEWDdgLxVJiQ+9UfT04L7/OItjs0iTx6i4dZul3qBk0wv
lpw2ag0Fly8pKznQSVFs9+mp6RUOSYmJnqg94vUPlehszj6iVonS82sGIgGYVhnokJ7pYbsRizEV
E+K3v7XrXM0WOAeFQeoFcMTnoR1tmzg43nn9Blpy/df+Hj3fN12xH7raXp/tU5jCDvR0lPPxeu2X
773u6eag0oszblIzJBLcL7mzteh+VCGKk/D3DEN128zQTZv/yIx1ePJXO0AfEQnnEOPEJebxd8A2
XbQFFOE+q4ZNnEspTVe4gOE+SSmidVG2RlJpAOUde1sAWYOyiGFUPdoSpGkJyWTcHxzQmygePZWc
kxpjFJ0N0g3UV2FsOGj4zfHzy119VzP8JZfg3LzFSHg8V+0zm3075dqCWyC+2ZMKjXK84Y7TocMc
yfXZ7y2j39JjKP0g/mqEiirdJpPQyR/esWbyloHhHZwXa118z04+e45zfsQjgLFlrTs7YwJsHHvK
bX7DzT/j1IUzWlCpZ1fdb9raUegotQwgo7cuv1nh5Sj2Q7k2vZvNTe76zblG3J+OxiCsP/bIb/GA
QHJYy1QXDpr7J9sX5fOKB9wz7md5o5LigxuHaCncKigfkJoLjejglrzwmpqt4EgrbNq77ALzVKZu
bWCSPwv2bS903lGmap3ymPtT43teXe5tNe0plCxKIXc0iJ2KbZVxN1h6/2b432e+Ha/lflYagqEE
/VwgoRnoSsMPGJ3qWWSwAbF5RZXozcHGdMccTsI+05Kr6HLYkuv7zan91o6RObjM4R97a00UTvNZ
wDCMgnpNIksZtSieoZdyfn8f4Wl9m2u7oBYp/88TVS0CJiCEshqM09LVke0eWGZgS/wDa25ACTk/
GEGuM+ngIhxMSfFcP4n+/pJTpW/eeTou706Sj+gU+uMa+ByNGhbDYZbMGeC6Cs2L5TiC+guhnHea
wwMpR6OGe92IFneXEZH6bu+2OcYx4XMS7DgDVyqJEf+uRzfs4NfDLfsg0bSJmJAU3bSUn3pro9fQ
u7ToNVaFpI7G9GYMX6zBHZyQJqQ6mjRCtzpUnCZSctc5l+weO2z4idQzFVP+ISqJxiZYp3QkGjH9
kBf1maiBY/sjJutSP2VJANdVkc1WCzX5JhwUm4N79/8GTYZ2YJzWfSAoBlv+R4P+x2WV4chlYEMu
Vg8ZOkyDyCsg8qulEh78ddLhyn3/4AsR8U4nM7YA2Q051rAItFA21r/MBntl9gWdp6iax70ssgsv
2CHOv+uUBgOrSj+OQx2zvRhh97rzJFZwR3ts2zEiTTQWKndGYMiu06OZNVnZiMReCTk1cOHYc2vA
rnzu8nI2i2DX9SgHwkrscrfi5XFGB3oTKM9sA9NBAsFL1XvETyGJtpvP4B+fIOCVX8jCVXQD+DEf
FkGrnYSqOkQ4I+VQcbkTDtEAJzcN2WLnUCFkZu3+8DLx7Bxl0mE5dHjjkEb6xnfZr9M6QpLWNIDR
4wGqBeOCpjlSi+chfuR3rTngCEqpk+W55pJKZrvHKuzOdETowS0JwXu1nqqZiJxmI+/VmogKyKJI
dbEhasI8nGDdgzrNdh1AG2HJWr3EbqJ/k5ukLsLnSa82snQXScv/xwgZAyU3yBOvqQcslPy4FrW0
VZBzAZHzPNoobLCv46S5aWq+PK8DmT0P8QZh4Q1ct4D2fyvBnVch3yne45uQaUSDlSZeOg9iwsY5
mIPvgNwkT+rDabciwg4dYpJyF7xnBG4Peqpq7R97H3w6fC1ow8q6lnTcoT1Ov3NJbKu2/VE/kfP9
d5XfJuObh9dA1sEfUrH6UWGTnJ1dq1BQweY5J+XjoiZlXWmHlUra11usQi+Wgg77dPJGmadEMZW8
yGsYFy5YJPETwm8RCaUc3VLb1TeWbS5IIYpJfUWebAHeba+XHVlbH/hRVNqCAOu5kRRGxrtTA4vi
8hoGJwdUIJ0iqVKConq2kg88DtIuCejXVIFyfN4xlGtIxgg3O5g+MFWVL/3YvFe9mTJ4c0+IO621
W7haeV1XS68g4IbQaUDRzfK1bAK0kjjc0vT9Ip5yc6fBXo2Tkht1slpqqpXmo7HQFgZwNnuHxZux
6eN+n0uzvRmJBn0ZNQqi4g7fpQteLQWmQ+7tRJV9I2NQNG/sCZp0HUtVmTUDlbRXr9LLeLePqSYj
0tBOgILPgMQeBGOkuX/fV48spwa0Qo46fY2hlkZO0Xv7v4QIw2NOVFCOokXtj4qXvophfMiPbX3t
HIufD7u/WuM6izUNJrcCew2SIpPM3xvOjzKNhyKq1AfMeqwCK8MIVLQhDLe0LhtAHQhcDMlWvicS
qQwI6I2F7rb2yx0N+fdbiKLeTao2TmcGs94VKSDaUQCFkRxYl2NGptcC14mcE2sF/5TBswiyzxwT
3MJkndZgWu3Wx8Sb2kR1k0pmrqNlrLfUvcJQC6cJyBkVdJsX/I7Kd8WUaxazuFKQiZ9CyxUZZ6Ly
73JeAIpUgFaU2af0y0RZYfmDAyWyz3VPAZ3RWCvk1DOz+9xXn/lNLKt6ihHexFoS7sPWjGYv96fA
NAoiB5cNmUOcg4xVr+M+ZPkbeQ/DYoKBe09dAzRnA8LVnsmKmTlp33kEDBojeIO+Nikj3/IzWyMb
r/Bh+LNUBWfmpMZlxF4FDuvii9SZx3yiFFs1HvfDnWc4nY6BTkZW6CXhYAeJO+0vS7cOazxa9tcZ
8pUkXo6C9Bp6lhOS2nVdvJqqvQZty4F1cGIozP9iUZk4F2l2sWyodu7835KsT8JRzBFkrbf155H2
yDwbfGfFdIrlevF6diw3fMk8pOjSP3256bL4NtiapNrzYrWcVa0uF6lriDINpKX7llWRnVVxcCk+
bSjQ5wuVSS0sIHSn0EWBQGdhi80UG/KfZxCyG+kHyJHTm+TKQGOqr8lBrQfILnpMFL+jgVKVRxvg
2t4Jdkbs+ic0g4AxhU21HcwfxN3Y23JlitFLi+8+a3Y51hhWj1r+gL5k+Sp0I/8EigFluatxppns
wWg7UqpkhIqFbpHS0T8vwCP7gXbaAGKldeNM5KTooXugB38a76+FN0HkB98sdyNeM7cavUxvBSbd
p5X509loPFEQDkLUU1cj5gzlZGwVK3SIFINHGSTpTD0roYQr8FcKfbBviqcwZ9Q2E9yn91Dby2yX
g84QZJJM6dWpUUoQWZ5f2eF25TAS6PzNO+vpJqY7lu39B9PKbRP1NYSyoxsmlrFZIoIQ5rd9v4Qi
VgY5MMNt2dgMbKiJhXS5QyitdboOLI1P0qsAtMyQwTdEObtbpYvdia/MsHZG39Il4h9domMG472Y
d5koF/lcrcX3COYe/Dxw9GpQNqk8xcpkd9Jn8NDaoqTh0r84uNndxTRnI7ZIEtdUTd/Jmg+Ger35
VrlcJuyvlyFSH2tPwez48PqDYSmQnQu5pzzNMqilTI3OTJh4YzT70+4Iq2TITHfN8M8R8I6gsM0/
NAmeu9QhC+VyuUAd+NwZGdrsFdNgp3UZRWsnwi/kBwLLPYaWmPqaeGHEgiQcnvQeNrA1rUdvFKVe
DBt2akQkmN+0fK3AKRfgyLaqzlmnGbrv1XztvGXGf17oq0bW8K/OVW8f6gt7DmwHlL7tUgG77QoX
EQT4UU19KcDiGeLY48fN/+oGoM/ghhuRDFbfnEWBykfMKerWxBRni0muGoHKOib/W1PqzldPddVP
MKUg1+/bCOwTJbUWTzSfu1SDd/4zO6R5rWXT7wRfETYxeN3Izw7x9N2FT5lbCcKK574FV4nbp4K/
ZpU/51GaX/iWit/LXlq+cguN+FV9FMDYC+07ftDKr31nG2w2o0by2EHxKy9gyGshCnMYw1fW2wVB
wbQVoKed5T+IgIp1jkEvCJFT3cRhYOGWSxt4qkGuvOUaFz7BxK3HSDn2QjtSBGSwC8hR0BsK34vc
i6ae4JNyU/GK6tjJA2w33Le+IAXk10K553JgkXQcVOFF9u6Bspi6ohnShWafP6mrRjmTIb6lI2oL
VXunQUqlW01L3lUKBmG14GJw3Rd6ywSHnMPbe9zAnKg4cBOR6CAmYD55ZbzkNQJ2RsnjhCXL8pHT
vPj0Ge5WGSEh3B4KtEaDo2Y2/cKpOuMqmlX/V2s0i/WsM0hdHFgsPsZEzGl2XXtx17dTtO8Vz/3a
w7y39rg5V7UK7T7cq1s0ta3ZPJkpFsbvQ9S14RS1ycfK3J0e7dM94Lx31gmY3opSODW6D/Zy6fCF
G8JVgeoeSoQYoFOzaMjeVb7eU3C8WzEXuYBP7XTuFLHUwPqHus5x7buBxPPiTlMT+GBwIQf8k7n5
IQTPzD0P44vT8v33XpocvDh7nXU9RpDoIPKNGj5WBZ4KNwso84rHWhuZgLGFLONY7OQ02huW/xbL
0onFkUdhdCcnZbY656DSmGeWQZgoq7GdjaHN1BLOndqA2sNyHtydK1Jwfope1AB67/6QZfW5yMQs
79hzYTSPpIejtfqSdTA8paxA52rATO8nPgZCx5Q3Kg5lHf9/Zt9nVz8e2tqEDsSDzitLm5+mrSsl
hvXG0XE5aidvtSrWA3N2b3ffHiq0SbHW+DIuB/5YqWfiqYee5z/OGVeTkFNmdmi0GC4j0/aJaXQn
UFJ+75SAeAg2oL7SMxBkvIwICR3KF1XtLFQHJWHEtwI3QqsXE7r9zEWZHqHGCZOvaxCsWZgakJYy
Vv/Yaj3OEFobET3eZATbFrJuhj0OdaUcPmyvNVWfIJaEdwMZ6YUAlO+ZybXXVzenrSKEYLRl64F5
i8GE3NZghErL030v1s5rMvZ0DGnxFhvgu3bbkLhtFPdQnMp8cahGCP3I4d5e/yuOwTB9eYcG1sQG
u49JFNd4M3gGlxL+mhs+eFz4C94e99AbDn+JRkBEBziAiIeUgQgYvGnZG+O6NhgK6R8b+EyXDYiD
CGbUHNQU17bVqdOpaN1T7uJ3CBVk4mgLCHl8qqwDTmZcJlh8T9zMtZNg3bUbP2xto/gMXc+E3HBM
BS0KYvZ0xU0AMQ92ogqPFSzTPWWsiwVySkdApeuzkXrQ5Y+xyQcS+B9eS52Ko3pZ4ykeHR1dGzIQ
IYLD9HNBbXubMOM1HKJ9fu5/8yVG94KET/Ypi9xvNAlP6gXjO6pCgWLXuj+UIDMbp/z7Q3My6VkY
YrgDX79qjDxAMEAzM6mR1K+hkoUR14wweGmNMtayw+BOaRvdme7Ah6ks1A2p+GJWsYPIZpdYMSYd
hD+POkz6jy5bXLSTcriPmPyTH2AtBdVYSflYXSINcuH1SWjZHwUvI24IT08rALXItRBYwufIVGrp
WODWCLtbRQancn+RalF+Ch5hS6K+HFEhRy57h+nz5jlWcO0ivcWIlE49NudWoLapsgGmOb72wkET
yHUeBODVp+5ySG6+hdFXGG281+JPXJjx15n/6P8G+BKxzzsjWSHbEwB1a3g1bwQNupgI2CilaCZx
kzSP5dw6bC61AOP8QBRGqSsUKcwHPW4EeLN9sKHXRLwuZCtak8NtjCf78j4HXibdOQf2+eOe8lbQ
hv3sRcmG4SpPDDHuJpvhT3LUQFgLzrDRAHwDQoOVQ2JHOBKLWxZbUuIl5s6DPoxITLMH+IYGFo5w
eK9BOgehqLdVAKUzt4esuzFITXDTbgT6TrYtrmmRs1RV24fc55S2uIAb1mSNttleD054ByFOXrzx
ugGdkBSQNdj4HyplK1hDJAuGyJFuYX0IVUB1yhIorI+2/2FKUcIjDTXHBNx3m+eSgk8YVYisfhp5
WVQVrD82bA+Oh/eWZa3ySHwZcVcDz4geeYLoLRSjywkZpksV4+Om60ocnrQUCg74jbht3WS3tSJ6
5/sYQJfT1g3TpxWRJyr7IZI4dKwWRZVYcqB7h/bEUO8alpVU4WDNjH+GReMkLp98I0ZgfRbNKsCh
7+N11ceBdbMOmTKtbFd0HwmaPeEomLRNk7UVBC1Qjc/FZKilqdemDTkwRL/Y12Ydg8VNGg/UjwZX
vK4AETIJJ05bKOWYK/DUhislV7wj1Y3dFo4u9KE08q/2ijgbtl9U2XzWqlKf2TGW6Q/a2o7SSWzQ
iIK6GGyTwzPNO737IZyoxL5te58DZehVzDj7HwNYDTm9yB7Nea1Bav0+goXTqLk5Fql4w5dLfLVi
fE/L2N5tf7OLJ0eD7G7aLTBLv+vCackQhidUgrBVBey/CDwcO6L+bTrJ5f0O+JrMCy8WyOYvSWch
HpSAdmPliHvGNMhmIvjYNmAnLovkIKrgnhw/MOs2lu27jUv0IFINYb84ZdGDDysEHVFiYW1atqe1
B8nPtnjTwAVKekAJOOP0vFTw5hHq0iP1bkJe57w3vMk+QUhrYnae51il0gv60yM+FqpYYfBvUB56
aOUtc9E51BzDljU0Gti9Znw4OTqYz50+B2/orlRIH7yCSN8qOEFu6VneH9FMzutEU0fRVW7hoRCB
1yipDgHVGl1CeIxIYVCJQfD2tUrwiED712biYxFs8I24C2swOb90IdEUuxLUHrF6pe7FnYgFHQK8
krJnP86uJ24TqTG8wNhD0Tlq7T9NxYabRYn+KX59f1Kx/gs5wV5elYIKsngBZZVG0S8Fiwa/KgKW
Ge4fGqtehQLA3l/HjSh/B0y5fzmQ67H5wJtlX5Em6qc7vZhEdYdNYUjoi3OSXmDi7ovH8462eLZl
0+h8xcmeaVh9sKyJEZF7bYRlZKhSYJmKuE5b8SEXSbLWXfnqs8IW5FIg1QUXFOnISBBNDEFWXn5Z
ChmCQ1Ni6bT/dIYe82x/rfeQwDj71Vq0T7mycSqEI2Y+vKLflDrhwZWsJyQkcSINUTn6WcW2p6jh
08XQXw69/BfaTZfnfHY/+T15dcIxm54w6TAlJ5eyZ6tUJ5jnu23NBHwslPFkb+loOt/KMhdtvRqI
4jzK87rxY7ZwiZJYlIwRJ5tG3ef3xT1T5RbcjkiZyBwy/SZD+A86JeKXESyUAdBsiq3Mj6wuQOJF
96KWuUETXr3bLSV1zykRkT4K9LdFKLShcuHMrtDhElpym8yqqkH/8cQmOAmQGwJNk7UQYrXWSNP2
dYXIp5nij5PPC0RGunWbFvz0Dxej776FDMWRYKb6uqn7NM2gCdGyWlKwBLrDfgZpFDzN65iK+K1w
bP8aJRerehyug2MAOeXpJtgbSWwhZR0q3lny7PcT930pvLzm/CPItZsmcYG6FuePAGplBbc0upeF
8wEK0gUBQM3BM4mpAOtQK6sMOyHfOhmjO1OXAzQ0mAnS4uO4U8x8H15KUG5mxkhwWnQFx5DOsi06
LB5/2DidMpyaUVtwEnqBxO6Nswwjh16EtlUslGgekh6UjofWfccjHBqD92BaVdwUw/LXEKh2bazn
S7vXRvjnENq1rOW3Rip3x5K/CYa/eNgDBIFC9S4jr3X2718PyAaicWdfJAK/CXSe7GVVO2a74gIu
L+U1cJBzTFbwgDWZaxVAgr7xe38GO2PeCj2qjzh55uwykIqKtH4nWObBUUbNFT6yG0yFu8YPKVjl
hEv4tM/3McSfz1aw5x7/1nJKYcDgcgORQXWjdAphyl3XfbbZY1Fj2FxIuJYe3CvSJSrc2xJ1ZFRD
xLy1gvf3jslDQiK0zx+DLG2RnnmpkzF47cPHdpZKjheEEaaxojZCmBcZamRJKoutDt1I+Y9tdCog
cw9QAX7RahXCylzg0ZCGx4HfMLA8Y5W6A+VedPzTEJpvnwQrSLWQ0jdclngHetzG1D6etbiRVT2L
DUM7jTM6L3hADmH3m+lTH8eGqekdTg290UVp2iW7FYQ7256DK+2M5emmvYZ2lSLpGW5nMfI5n2u1
uPHQipB1VV+TChvax+Dt3bkTq8ZUbplSBfXW6/IoAF2tuukM4mXHP4MoCmlnOAYhmKo12p4qbdlb
4g8m9vORLWI8HbqHJMuWV8pvNjSnKrtG+zQRhMzvIcdE8lE2fHmqCa/kcXJTCzg5e//SMJ6xAe7m
S/8gCBRLFtxfS5yDcIHSpQhkpZLmt+/LnPztHA9uWdCIEENz+DfGmsY0azA4QFRkFWV8cFuoyCyH
3EyJB9qFsB+Zbhx2jqTBr7lWgd9RBVNMvVXNIfG9/ZgH/nXheTD6Q9LXt5RU6N3u8mPovMKYbUzH
jbD3sPxL+FvXj0nMS3oeklV0g7361RtU9PC5D+10wBInkMiJw0W82EKwZS1yCQ+fdQpWL5YJWth3
Joj4GUJpsGv+fGFLc/c4RIxaTGJiELG9KGGZ3Tm1+BThL3Ib/mwwBwlhif95xYBaG2SH6RNJqF9Z
dK5GuIEGAVbi5ckmIxE5n3hrEA4ggPAF5LhH7EUv7NyBk8LzEs06PurA15LE9p7JK5J1/Y9zg7Si
8LJs/n2LJAwqktKaXsuxeSS7UXmDZzQzVtFz/WGy4OTiqoqITnaSmKS18CUmF68qkal+MYi9oeaz
lZXjCwKguXJimTD367+C4FiiFnteoQCfeLKaP76eJrQ6n1vQCRRnMBmzUMoqCvk0Cs4tMbCEOSQD
IHyi/zIca4TJQd5LIxHdKATmwFQbPdfDrVRbb4vnzevfOVTfp4g/F4F2ZZbPvIMXteFnE4i98iQA
NqZm77Su6/B4TJgHgtBJ5UXlF3wKIrH+BFr0lWQWLRjrcjp4cf2p234jAovGn1DaHYeaM/01iL0N
sBlnH//pYTWJybrURKQhfiSdG9jbrBh3UaUNahwjD4smwwJatOA1RRfU7U3/ihf1dESDCpjdFX3q
HojVqmp45rAgzbEMYzQj2hsB1mfoQDxtTvm8qTkedONJJ3dIpnwd5z7jHkWQM10DEvQGNHrNyOHQ
QVDtekKpcyuTutvlD/7XUkvpJew4vn9bIu4lofgsROihSbbkNypwznXH/yZBsc3S7GWlqCJLZurb
Sr7dQ+/xyMPidevywPA+ZfjiZahx/691pzQuvuFLByApZkoEF7bC8KXYS0uHXZtIvpiyUcev0Rbi
VEK/QFex1ewGFZzCFcIF3FAp/LBIzoNMvkuKtzv1xJTUX/hEGjbCjm+NOWzQwGZnerJxoGGxjCmi
9Ype64nbGdqW3sECXESqldwPYxZ4lXX2pHyWhNvCxU4wGiJ5Y9//9ObnhE37pzLdvloYRKJbXQFq
ey6xY7x2CQYnRR982nAu4B4M5av5r/f3yCHng2oIL80zx3JhIVWqhbIpeP25Ei6G5pG8NJ94XUQO
RLG0/AtIpOcw0eioj835uMIOHiiniNxkMS0sj/586K7CyGWi/DQtHclrXeN7ySAuqRNTGokBEcef
IqBMRNu1vlboG/AN/4vfLM5IuCY1r62BsbLMONzqU8zprhj5iZW4wX5zM51/G2qt83Yor0rgUOEK
Twv4kowFZLunnOWlun8QJ8iNRHFzXENzCfkuWffCbxI1aGO9QpqgmH2ynN7DDVYKP15snya/KBp6
v7AMiJh9YkLq0ibeYcIiNSCLY6BIuwDs/k7Kk74Jd4B1/0MyYDAsWBj83TDl6QD6v50FXZUenFEI
EeH+ZvOsjNxNrHw02vYoCoDhB4NOKKpJKRJkl8gkNILZSPoAKm/OnC5pr7XdhaOFDWmclh2+q6xA
uzjG/1oWzH9sIqfYf7zh8j5RHMco5RbvPOGZT8z/RHNJxl6GV41UZP/bUHB43ohHtHykGdS4LtLd
97UwfN15U6UisvNG5D5IFBuCK+7Ip72PiN5BmvE2RxrNtkG9HaPP7TSfCOW46LheqbTd66B6funO
icdzBEkEJRm/nNzJHOwqZ+HsW6bEVFtO/AZx7gl5Ree4IYR50ys6GmZiICdL+Id4JqGEjmdiKi+y
3t9nlp6X7Y4Phkb2pS4w4q6uSphUcO0xqxFp4DaTrzQeqSxwudZYxlZmtJrC47G3UMQpTlDaVGbB
HU8xhA1kM5N9tqGEuDfr7y/xQgoaBnLTCoNoC+tuxIIxIfu/XTFoAijaNBx4gpFvpw3Wzg680fl8
Y25xw2YhT5T1nY+bfBhdsz2u5bMeZdmxqqhVI1uTBKHFEN55nfXIbGtt4LJ16EnmlX9HlLSEZu0E
4bu0f/NkM0dbORi2BXoW3Bf6yzTQJcx/5cV243yHhTKfMfTABOGakhI7aZX4vqUKN/6JtC59Eq5O
rXgW6xLUA7iy9533t2MYM9OVF8cT/Yi1/JpAMmTfR8Y928fitNYYhG56O4VZeDiIZoQ6Jc9c3lFS
bwBI+SxPR1rsXQkEdGJ0MD9JFtbnyuxNPJ7WixTT/BmeiDJO/87zdzDcWj2oik2s3Tb5YaFbz6IW
4dj56LraN277C59cNGEck2gTXsxrVCoaOvfPaW/7tuOf/q+I6bcrfjuRc6a1orM55L9PCvwzXLIi
V/n5zVrgvEvvkv1H37JMuyBASimuo2DPlcrBZdyOy4iVMiPHTS23TZR1HMdSIGQbgT8sc4yJEgOZ
wOpJy83rD5D5Lb13O1jqwfFFzJkNQLVkN8tSLIusYHWsgp+dW3TeP7+ihQJFcam4Yv2ZG3xHLIUG
CZ1kSAEtHhkLV/7zlgKenixJyA8o22G7m0rAf4/6FhHE1m7Yj+DLW00JbNj9LR/Qs/80AtpoCnLV
oFHGdhowWIvXR8hhHKEKV0RL3bfbSNqg9LSVW+dDzCfhVmPCUYNh5UL/bTIrOMg4iczJ09P0AA9X
VT1Cb8aeeuseVIn9yMuz6APNh4xkLkRyM9EWhcBdVrK5tGo0CCuXA0A3DCh8e4fwPJrpq626OvSP
TCaOUm6dMBjnvrCeGNU03I5U1pqEbrU0GMLU1o7cuLJWXrQsbyTl6r2RwpQtvkAT0k+VQ2qqikLc
i+e/7fxbaiA6oNF1Lw3a2ilpeZfp8dWDGEF+fdO4u+aElKnnYD74SGXfVdBZWsd9nXvm8KV1a9Az
LXXgU6rYJkP3jQCT7j+T7k670YtFb3ls9yFsX+4hPMcF/lj9JT/gGY1XDWsPlYMt7lSCTbw6VX7J
+1tMh0u0HvUYlVzXdwiRItvg62MIAz2N6sXJ1djUaRFKjfvukxNH5ko/RIKKGmoZUWh89aWsnI4t
qU9m6EPfNoc+06yE/dkkQ5YszrlGmrUBTHyMuIQA9jXMCINi9juKz68FHJbDSSqfSUW3IJnOGVoj
glhx/KMm7klINyR1A7d9B430vAG1Oy7Dhfqzzo8PUBJjQkuUNzHO97qI65oCC2c8TrFvNn6lXy/T
nMZmIbSG43+x/NhezM++p7tXLG4L2CI51Hsz9j/QDL8ZxGTzcFWQt9Pq5Lhd0OoJ+GhdqtB3MGO3
KB+U1VSUJLPVXNVkhldMTKZFgnAeAhmyBgsdf55Mk8gP+eTu94HiiQ40X+FDkBwM8qPaBCW55k53
Vd2EilQx30aVlh3WB7EuEabWf0kw071ullta/DEzU1s8LaKCDTkc62dKhXQlvZzEndGI6ClznChv
g1Nv9TIYuYK4C2oNONAGHg2z7SfoEI5N0iM80CuMj5+7t4j+0/PGPy+6Y1Cu1HOk0yDBBf22ugsd
oaeilpzlYvL4Ry/PM2stnMVkpU1ZhPt8SWztjB3jW//wqnQfijzClulAyu/Qxc5/WPSuLABM0HZ8
/v7L0IX80rdGAqbS/hvv/vYwxQ9r2TmJSRBu9HC/keARjVkBEAVzbvtbtHUPX8Po5Cxt70DsB6V/
DLjbsAcrCEoE4VL+46MDXbxZHoQ2iSWpwYTpMTRmnN4ix5QS3K3XhVL9FlnYmoAoKozwgNCMwaoV
gWGZ+zNIZOb/5b6pr8WsuzNvwb4AcS0FT/EfUlIebrEfBsZNnn+uSBVIsfO9+BZPs//JnylpWuhb
JUU11tCot5q/72cGfT2I1DlVbZ8JsR7NGmEqMgBMnDg6Y+MsyuErSngigELEQSELkmt32mXwE/Oz
RCwwmWHMY2M5QLZ2mX80UnD4HUA8J7wxR3/XeHT5tuBrDjE0MWAYcxDp7+RXMKhWRsAmk66i78t5
fLSY8jmrfjsEqKfxx14I1QbPr1hR67k8NrPqpzKJNeEjem3Exj4UeOfgv0ZdbOWRVhrkDfKxX+nr
lBeYxbZLghtXK2jOMUSYh5/5dodOuhPNLba5b6V7einsC/g7aq/pMp0kEtzxK8FB77hyGXxgYzax
kfx03s+IVlF2wU5CDK87l7m+KZizVphqJ7R+Mr2/VJjl56PReh3spXz+WooJh2eVw+byVMzvlIpH
cINysYNLuNB+H/G1ZQ5rtnJSfkmE1tLnxLHAiZxThaY5he/+3VJYvK5CgtylIkeGMR6rwTvVwcRX
aroQrbkNi/dTaOWQm1SzMYGUZC/QHTjhR2VgZT+Mqlu7kBRwi4e77+doLYgcr8VDKI2RgCwWA5nv
pLHr03Dg3e//p57kNrGlD/2sr0vszfy1AHcifFyaRb6HE0fk8Msk5JZ+dzELW3uXZZoOQPgnFHGq
YOxrD4fSSIwCA51Lp6pu5td21k/GUyeDQtlDHHXB+VIxY7laRJ8T41P6BPCxhRuBt9H76Y4rd2QD
7NfMubBlBw7TCNN4o8MSRwUVWl+dnpJFS8KKMiHhgMo+pBfGMRwgK9mAy6At23QwnLZGbv7spMqL
Qztt74wFUOQzLHp073tDOGESSeP+N5vdYAsOR0QToaHbzHvgbc6ngymkhma/PfuIoUAFRKLRZWsB
UxDmpYMYsJY6nVo9vtAdUkzR/AMspmBpYoKtbzCDst9K9JaATjnAe/VsLXnp/oRRC1BTqzAaNG5H
fj4Sv2Vfsp0hLl7O1AgBbMQp41kf48QcTn+pwDAQ5AO6852yxUrYeNGUTXSCyw/8Hsa1/TsBxa/O
CMsMfAqORdjWj3TUBMaUbDcScWVai89O8rosd/ds3GK0pTG458RJqfO74r+uwmMBC2UEN2oEZJ+T
FnDE1v+43eRWd6+NLZgIItOL+h9q4w7wyTk5T/rgDv9BP/a2kLclzNPFPf7I3KDBRZhVidG9oPr7
ye4BjLd/oOH7Xuts7yMYppb0Mh/rCXGYb+Z3p2PJ2t2Op+qmmHz11onAkTrkinOkZyx9BEltptEp
Zjb+w2ml54zl6x5u0UzwcqukhckoXlMW1hOSJb0l8beRlUzR50YjjfLbtbXgVetORHv9Z7wx/31D
z4ooBN3s2eEIBU2JfkrFjGK3cP4RR9xaaGJMakn4P1pOglyfZTWYbJq0jiivqAC9fu4OqAqk93o5
nAcgMhzv4ihEzBhS6IjQutJwfZdLOeC/QThFS2YXN7c5COu0x+VwlshG9NWFQqiFctSyu1AA8Vm4
DUBPVF47hQSqjOFKsbWCo4J1tDoktfWkj5fQbAL7CDQdn14EFCT1lSVtdSWJK5p4/wwDSxkusKfy
GveT+gw4qR7WLfgN/4L9Y/dIExnhN8sbnCGbloWEQv20BKRtgS0bTUOx8WCuchsC1ZaobuSyIrLN
Exde6oEsGl7cZ1t49ulwgSNxWXhuocS9h2cc6cNZH0iqFOxWAyzi/jTC0uczQOrx8sGo1DkJ098d
6rDvHnG+xdYoq6DmI3KEw+6rl88RO6b3CaZsIwkbCtt1OF8YN74gWYD6ZfUAywPcMIw+LVpLJOXS
IT7i36d8xR5bbGIUlL8yfHFxYciUEBjpanUfovDzaS4GQwo3X3Ya5+4Sn0bDHzkrYbYZcrOsl3/2
VowFPneFw/GHoPJqfDbSVAifs08yrdNE25MRTfO7VLB/sDe16bBSHBrloTpgs+rt/ApfPzk/fUjY
L+DWxsQy9l0rfiCCo6hbG7Izc+QJmXzmQLicAv88kyEa6LV7BNFvH6mW+cSY/k5e4Jy/bcJUK0db
1SsiF/8ZJpd47UsM6C7JQwfWf6mLtD1FMeyv2noPFlKdVQ/DC19TiuMNxfnPZeolDBfJiqKeyb8y
S0UpHI2dkNagA8JX+7+P+iFJeY6Sy4wprT/OTKS7D6yms8OmdRRyrVj2FdbyGaL7ShNZsRJueZCH
USsDifVPCZn+dMDlYQjxQiYcuplQA0EWgaqxnJJdvPbV0CpXIZYDlQ/UAgzMkpgqwhfNIwlJnbEA
vJAQnihx/CmoPsnKkd1r/AM+V+2wbZs08cyT+qMZcmM8ApbTXIpf5E4txZuEr1AlI9wNnhH1Eg1O
2ccve3xUC5HVSqBnmaZvkKlf8h3eAcrGqPi8OfyX6LFS5hr6bZuS/L08/01GcdzOrGKS+WNTQhc9
97k/1iu/QYUrVWePbAJ71zpJdTY8yFQLF6ioOdvGOiqttuMJIgNSLsHlfDXfu9+7t2e8TZ6MvQph
ndvlHxCG12rnD+UKg8G4uS85ewuQkXX1/R2VlJzjVmVzkPvc/0+KhKkZjGEddjCoVh8SKJJhNsK7
Zn/Z7qf8CLMh1Zf7A3KOd4eyabxu55lalzYSASBd4KPWcZclg7mGfKW4WKfWJK1Vl8FH9U+pc1pp
i9pfIrOclIkvotfcJ5ou1wK+Ezm71fskukjxXRjeSJWeV4kMhG3rNiwylaepB4lYZxSLhN/3nedK
5TFy05NboowVkU4hsOq00ERRO+3+dyqqh0cznXtjd8MQ5WWn99kVl26u8vXRsnZtIo6II1g7yaCW
9uUofYbZA0jhqpNMMqfmEdwXKXL1DamCaGxvQXE5JxteyzSwTl5b1lqgVB3aij8k9e/Uqmteuc6L
HEtfIjFh1ngMr6GlWoa7/nrktwGNQl0uG++wQM1sRxb8aSsZrfUqya99paUBNtha/j/owAnfa3Cr
lkzPLjh5BXgl/szU0Jzspp0ZZ47B83x4TuVK3YrkvH4Sec86xpVy3eYrua99PrTC1FKG6U/1/nhS
DAioEhz8/z+IhEAfMnpAvlqP+Yp0mgccFdmFys3N4TMzrGp4ZcVm+KE1lbeDXbpN78mb3o9Afbdv
VTtsgdOm4uL45gqQVmpjnMLk82iPI4stwpuEvqL5Gm//A26aG7EkPUtG/CS+iWheRDP91vszwcKs
lgFMRfFkMxuPzTNhFrh1VQ9UfBDlgV0u7mDs1KS/STg1cznn7m58mCU4d6BkJ/PNLjDpXRY3W5f/
nvcDmLDo2waCptfVXgSpO2suBj67y8syTIrkxc8L33JBaRNIDjB0/2qYeyqQuXow2uYo9ksel7Rn
I2Fk8EOIP894soi1c+ia/9DjqJvY1e16RXU46yjAX0sDaQXheY3j3lrTR6+mRRuzoYgDFij/Ngoc
b/uGAF+XKqz29xF1nT11h4xtBi7Oo7eQgZb4rFRyDM9iTMCEyPeCDi2XiDPH/kmNMgQT+usC4jt0
G1JMLNbdjFxJuk/FrfyUEFDCYY6YBGXMT5dB1H+QtG8bnM6tVccfBcb1EIK1mS36c3RNcQ4yG7Wy
wxQh4Rrzju0HzTUUFZt/9cRGkxk7UA6hph91czsDOyaigDQFWbs6+QVSJwqAQLKZwpGjtl5yezDU
LVmnrOhzXsV1G68jp71F57Xby4dN4J+5MHPm/dgbDzXYi9cZcoxK4H1u7INPJrn5rrth1Iu9BHIK
E41Vscojxvwfxw/s+n9X1FeRttEydiQzR06k1M03YfW20pnjhm7RFPIIuHMEA+Ip4hExb98S3muZ
yRE+/JKbAJIrrvBysdhHoM+cZW8osJcgsb7dm6MGMyGvcb5+3T9BAtLv/GdQnPlH1YaZw9wtFNW+
eP/HmITmn4yU6ue6ikAQyqZs6RrSMA8wvZywU6MM9JS5ZIwwAYpmcM6eFT4TrDntb7OaJDcJcVl/
9y4KlsXf1Gfmasj4kbEI8PBE921CmmeubvKxboiEkEZxaqIYIpu1TEfwb94stYhQyhj+CixH/DmD
Av+kSTLzNx7gD7dp7eM2G7ujxRcUO7NENq2OANFNYeEysq9qP8icFPGoNnZrKny+QU3zA0Dfq2x8
uy3p32yTd3XjEHKNOBoWC+qlB8oX5vgwYcmHN/YO65wbtfwqrf1ZUWV2FscHzC1fvTwGgHqg6DU+
+X/P8+wdoUh7kj+IJUDaYoXDdyPWC9bCKORU9dBK5Wo63Y3+0goBX5xz88h9UTDT5hs0xSboepmE
aJpaERJJstbeNtPeae7BlqYhWOpT9cK+ZlQ5DKxS4UjrnRBoqafBlS0Fw/vLuEvy7VxBdrJ704ni
0iwiTB7g4V7cToeJny0pJCBzSAfJD6Wjnl14ho1zcKgjXdA5KIA4a/+HqV4/VYxclsVlqXo2W3By
Cj+mGOFDFMRB/r6TC4QyRAvmOzHl/cxbbrY1feAHnKVnviaIa4KbmL2dOpYMhrV9BCIjnmihGmeO
nvaXSSlgPJav13GRByKLJfnfd9S2auBm37riqTsKP3QZaDA/2vzoubPmG4k7Z9g7hjQmcEMGpv8C
PWnm5WSUJZ/jWsncp8x02WPqYtAf+7d2nhF5SM4Qo8BLBW5FGEMotM4uFxR7QWNTuJEsJgEAxv/k
MpgKz6YiSo6hwDiIJd+d5qX6CdcIyhGGKPVuo3RSEVvQwKWKSzP985tnLvwmi8zJznj/DyQ2FjYB
LR8rhLFgFYKuPCVcrpRDv6pYx2fQvd8xjEbJ3mwV/08oCS3rxSfgLvPA3iac7iIe+5FV9zKOo7Dh
WyWrZmRIrifl+2w1OrkOoWFbFLJdR7Ifs8urGKhiNAGfGNa7NJxBT+FKxQI8oJscw1X32jBh1Xvj
r1q1SlIznzaQGxTOLDHnY6dCBJWyuwYbwWUdIfEtli3S8af6tZhx5jzNY+l06ROEyXHfld+6jsPU
0vzab7s8MOOylw97QZMMaw5zRRZVR4MfiHYkpHU7vmGbH4HnF8Y6FB3IqrhmzD0Ldvl/PXn8vvN4
JfgA6XzMJw0Zv6Emz4qn0lEg68Shz1ogDFnkPsyagbBOMVeFYXSqo5GrmMnUzgEgFwf75TAhxKZ7
IkL2hQnH/PJ9MHlGijMlJoSdNg1xbokFCeJ6Yqw8nUIfEOyg90Co3pcvHUf4NLJQW993I36V5WyG
gV9bhjcr8XJgj9YpNfvomNHvTson5zOp3HHQPubiNAW4wNAxtZdL0CdOz0abWx5gfEW9VX2QZITV
kZOKxfRgLKBQtnNvpYSv0EubslduB/QD8LROTh8IKI4AQA3TN3hjr8yr/8h8aRqaAydNzA4ndq7J
bGVVs/TqFz0uEUEUA/MIsk9jwK/9x6VulNOboYgBQQdIr239TjGs+oF3vLTvGQKekDsY8jvGdzL1
ZjYybZMcvfk7CN68qKjSZ/EOI5Acz0vyzkoNWQ5rGdtQUrV7wgQSLwUqEdrz0d6hCI6fldOA34bD
yX6He5JR7hN7WTGEQIAyYTi/wDofW3WSyvhnlAW7BjveCJKekYeW/N2IMxVMSzs0QcE4p6Z2iUWv
ivrmR0XNBM4A18Q4MkLsQWbNJ4nzvXHYQADhlKCKc1BeCSuPMSunzye1hymR5mi7bfcxzl0BZcnF
OJenv8H63Xt0VsqJOJTEIanLtUbI4XwMAhBrJ2Bkq6ZvO2dHCzra7/eot+D9DXKtBL+3QPKFTlb6
SzZzGeEvytFhQwd3QFKae2VHIHBS9G2aFCConeRd3M6SEKKddgvaHCEIGDIxCcyWbgTFzHcR3/41
CLSln2DpKWaGvI+ohVXvlprFK4DYsE+luReAcRnjMv/40tOykLRYeGsZtlQA3OXUFGdL7ajIdLiw
XLEaGRy+40AXVEpBxw9As9JZqyiJZw0ZXCLNa+Wf/bKLK4EAkZu0PE4gziAQt8XLRk+2Xvm7CHaL
A1lKjihxQCl9KsTx+zBdOJ+FTjESnankH1oDq3q4wb2vVsrmPoiaunYeUuREmwdGaO5KhpDYlcPH
yhfl2Tdi2Ca1glGBFxyeKYVZox8USKv6GyY24g87L+m+O1TR7+ms+FCMg+5iCLPJx/Bw0phwfr+g
UeSjQNnvJVK5HryKmsz4DlYWrbgG9kGiVIxzcdvEz+5DybrH6WC0XcP+wCEI6FL+hcG9G5KLM29g
xmGYnPIAEc6o3AfAfokqHTmDo03WCWbwje8DzoRdgWkHPu+fqoHbvrr+SON3bHWbZ0iUc0XZixSz
qIT8Fv9n6kmNLJc4CKKIxmFQK9H1wD30ykjalptbKgLTw2jhMsl2MPhr06Ao4TSsckvCsY2My4OL
ZIgszoOn2WRY6XsOa5wevYCY28L83lTROFVueXL7QNBTCTimm+idWpHzrYg8W6uS3fXmIWZAcDry
rjBVLNAqBIcHTk3zFa5rB6ppKi3XFWMdp5ismhc2zp29oHQIJsFTmDd2IsQamKDQjk+PIaUw+05m
iCY1I3al0/8qG+eaXgekcBNqMKArzc/ttKMB8JbEcCrSPADSxyIx004bUsJ0468O5F9fa+AbF1dD
1Aen/NSJYA3Gvg3l7NQMdJH1AZ305l5hnvT05MsSrEmfI7xDtmFNmFvdqyJkOx0644KGF9rvPbrQ
KDRGtW80iTASYLqZDBZfDzoX1FuZ2M2iMeW7/Vfxv3zcxiGIWtEdAo8cmNFiV9X4C3XsDTJ75+2D
25HoqZQPye4Z1kRa5w/W00KC9+pr0FoKMgZje0LVbZhWnlnC4qWVa8SKVVfNUypZx5MmB0sM0GPu
PDqPzKO8G3LXeXkGMYUflblmR1TeQ5rwf5GtFIGm0AN9/QdJ4ZYIqeGQOEAR8rvLdRTQPP0JOsLQ
iuYmd07ncALqKEKaBR6GvwMnfqU1xWCRNsM8f/A5wi3kTQGpjTb7Q7QMqzdkxElBCB58FZbDC200
YqWzAi66bI2ANLzoUuDMKdVMQMfV7PpHTGUbIidtbn1IScORhc+XdrUmWNdqatLm9SIGaQt6LJLs
CFZdr3Q1bBku3BaSV3A4JZQVdJwfaJqZiSdZNpRjoUMnm1gcXWL1lKpM+R/XqAj2wjfXZvAC3qQx
5sYO3XPCWzFO0sIzXM+0Ywn3TixTtomiwJYcm1HnDKOPSKOsciAgNutwIAOlthI3uePKH2hOqHg+
PBn7QdBHTA3Gc5n/kyLZxYAEwZ/5Ig+Tfr86d12aq9UNA3KI2o2fy9UsyjELPxY904VsZC2KkIeV
sw9yBdT36q9PIGx2f45Kd87YdBSTSBaNurDVmyMQ9Cik6TnpWvbPc8pZPitIvtbDPXt9/xdtiSNw
Lg8nceLl60y/fohCUx69bSH3jVdCRLnfpaLAxS3NHChtygJ5MvccvXOWx3Z/JQk+nZa8t85sObB9
7RuUrWXzUmE75ODDhDp6pjAJL43d6T10eIyhD/cUaK/bg7b7AuOoeOdVCXe5QcGfy9zJ1wrh07R8
M8qnmqohVcIAGz2dQI+n32OkzhL/nruHkrs9td7EWpTLMvc5RaapMnpEi+A+9e2gz8yM4L1gWs9q
CnWjaciFEBy9zd/31uUp1T6Z81ZJSTOJp6WPI9Hww/hClNt7kL/YuQ8wGuor4ywccH239VJGIGPA
gravNX0SpW5+LiCdD2oUuzaH00OhIlAyokrhVu965JvewOS2dRB0fyKM/t1ijnRLJI1yH2eYQ6Qn
nYt6aixZYJyWjUEZcgSpfL/878bPHB1BPQST3pzUQpIHpMt2VQyQyo17EYbBotHPWxm3PGuwedtD
8g09wyivCzCw7EUuG1MSjpeicZ5DeV1uS7zyKckGDTHr7vEo428RMCjTe9OddfufbcwO3paarhCn
URfqVnXYnA9J7EHjclDEDWHDvbC3G8hPyaH5pyHSv5pvfX946GRONZI03TwhvAOzMmjubtZNRWf+
FwwZ+bg35hHm0GGHfb6yfEVWQUfnvfoI9yGhN1svGt+G8sHenF7BLdnvZliifp6mz6fiaObb87jY
dX26VXI8UaAV5SAMZdqRMlqhEWW4h4RUsd/PZDu/bIkkye48YK25YCkS9SmG+/sJIoH4ORwcklIx
QWeL7PW6cy6GO3wLljiEQ78u3EJ9GQVql7z11tGgKsmKA0Me5DBGcYcKjORwuINW/VKheWLuSx0+
rg4sgsUjFh1bOQsrH6MWmoBImSOlK49VuXWPCe4WwO20Rqza7CMcdMN1HtVp731c2Y2w+9XGSKvO
IhGcwGUaGGG6T9uFmxGjzRFOWPrYVsGCpGULkKLwzvUufGsjuVmMiXzT2+CdQYj0OXjkQipj13me
YhOHpQT8RiJTukJCsxiI2xHniUY+wXcea1mJ2RLhk44sKYWqIwTms/iMQgz0asFsr1Zb84nqiPwD
r6hCKHw/L5dHtmsMPChR9BA5CBewlpuariDIgOB/9HE0GR8AJqRGaEeMs6U2Uk6T8Dr1ysvoeP81
pP3vjPRTTO5x9XgcHenBeHUcKSw7DcyIFeJdhAwDO9ohf2OYx649cMr/3DgCmhQPnBxpvWdwh91d
bwztgUIKO1ohkW9HSEr99xsBeJz2dP34AcOpSGuQBETrf3xY2NDY7Cv5Nxi0g/sfEB87jbRHTkWa
X1uyZNt9FBZlqyHSqhlO9cEpalRd2/hsdEfTAGwOL41iwSuJdio2KOhibZwAwmb+I0mXOpKTekNY
IpuVtkXMj5pFEhEQi5D+1PTyuZji9jBxGyn2q1YKfFCPcE2R5vPZ0NkThRR2mTgBc2cm+dsHd8L7
8W2ANwmN6XsOZM04A327Cd6koIVrynBa2sNuIqC2TJ9zvWqsGJtnGhXrA6drdLiSIb6pB2w9ijvo
zRFKRF4GPRrZqlwiOmVBvlZDQTX3XCCyhcP9REeYOnaT3QnRAqlHElX2JsNaZIyzkCrGtdg2LdAd
Jr0EOWrkUc2vHW8sv0TthqMT9zZcGFeEAH4EkSbush7oyUHV5HINLMNSSjGvCxy63vmBe4iqrY7a
yhU33614W20CEMyciUPCeBJFqerYDej1umGmQR+gyCgQrGQCwTxg6TtNVoqg6zKwIQGSEYdh3UmK
1ZhN1udkW8wZKgHDAqWanFkb+0DL449OlKAirTANWwOH6oqOLBtzg8+K5OdkRNMxv8vrRY6AHpUV
e+PxxttqYVvb7mdkuu4PQAQtigfgRKZHz2lmctWerifc3ox39giQvkp0EEEAKK5BQEsgRPZLbR8w
3hT/bt9htXcau9WjLir5COEk/JJlvBDKGRqIDbV3isx+tv75CNwZuFYIns28K7aeu5HN2e7yUNXX
CLfbwYDBik1TKdYH8xiOmXpiw6QZ0TpkoFYdvsDS3L10FF8QYVXWFZ9qTOyMo1i2NI+2Q+lWVSjQ
o6y3qBl1B5ng+71kAjuoTXjfIPjZK93+XerDqvR/2xylHDdsBnS71ls1LkEVJ/ShrR6Mb4tZvL3n
xX9XVPC0z+HWegIFoWvDpZ0VOPQ0cJ6LHEUgpf+fv5AJ8vAuafVLINCBwDI7AWKoEIqINqWf5U4S
apfWTl9RWx3HnL2paX7bOYGH8CiDqbBr4yAROlL2Mh61flY5jdc8D5OYpaBYRRxkvMUOAjZ0GOWO
iEK2GBKgRDDdZsD0NOVpGZj9vZrFHhOk2CwGaaogO7MAdxQpXqnCk4Txk6Nq3+tFeASE5QGyIYCP
La7hpS7Wo/tKxfwYsffKnQrfqzyjVli15/LHHcmzupRbhlS9nDFMiG5sH07JkBvW8yR9FLHGHK/U
3O1cy143lHXVLlwp5l7nQ+4fHt5yfPWDxBoCo1BfMxbuTv8aaMZx154AYjMOCIXuRDeeDaR4BFKu
M/UXOEHV59U58Sx+RImvazRIQsnyfS/peo4vwW/pMvKR0fRsT+KzU6blog0n8sobd+Ae5jdcZw1L
ejt7hrxVRYjAw/YbJNsJZZXdBPooAn9ri0jGyad8bZ5qyng0ijkQ6Fwb/oU00A11SoAzWXIf1HzP
yoiG6fZs9Ef35N1uF+XquCLW8OjlCpsbtCNmREZIE0lkvmzTDymz8LEk1wN4em74lw5ig1GySmAj
fHdXlWj2Zok/+9UzmMYLbCmY80jXKdEoDp7p39lXNNjt0QSrCLKc8fyxDYVaAuFMJLhnBonK19jf
zBNgo9ZJmuNmu6yBcyvSHELt9y0s0pNONO+yPw18MmnN6oWfRYlGTMjszTOgNnx+I2le01hf+hNK
7xJjd4DZRi8ePG6U2HTGkgdw4R30TTIJfR2E4Ztu8RPMnOMiuD0eyG2UnUcNIjOBZHnBOFqS9g1r
/uqlKzQVyRSzPF391bCk8QKkrFz65UYphIj3dKMpvgQfg988qTki9Zqoc0lg9yxCpmb0V2DWJNeZ
uUuEpTGcu+Sgf6ap5oVTwtDih3jHskggFLfhJ7IWeXHxH80wz7BYuhLsbaWi9n15FQD49zj+2MvC
wKb9RWshIvrq+RtyvDZJv3WIcW2NHPPJ1UUay7g6j/ygu9Ump8psz6dCl7FGz3LQa0aWfUOX0xzy
2vcyZ5bx7nk52ZgRAOhNV54HqqCBoH8XszcAbydEwyscF+54EXduUgb4j7sOgOQSvsjo8PwA/o+x
eNsc7zOZsOhodOiuh8YU0nAXj+hdfFMs1IsaaqvoeElPD5jMoGEhE1jmEHltBhaqJ4LRLKMJaqpI
y1RKN9OOFSGom72giLUVzcGhLbqvsLXFa+BuGF5eHS5cvwGRqCpHr78hurigt7F2gpMRpn0n3LGF
OoTBIkdo/WyIuqX2MIC/TtQaDm4JGPjyTzVXdDORECAy32qLQWmv4zInAtWMEHxHjQWaFWo1xWTP
7QzJPqqZzgwk0WYdecv7SzEg813chkaLrK+Wbb/hAQqNRsPFmMSETCa/WT3mzIjKv4mP+kTh6HVt
7Ke+sXog8H8jgADZELChM5Ya56UouSHFfM7/uoBV5zBvW3xsFo6bVWN6hi9N/Dw/0cD1SIoCzVR1
Gmcv59FF7mIX4Pis70eA1DIGvMAX/WmfJaS+sk7OT12wIJyciyMYvXbokUDrRgk1QKsx31mHvcHd
NRMDYQNTIrDlTysCsiFM2QEFg5oaiQklAS8lZk1KLgKuaXVsqrq7wBBehW9HH/40AKa6bZ1/7TJw
ZXWOXHZm1XpidINuqRGWSjyR113YZVrMXFgRmWwEhgIQbfXrsgM5Ahvls5wSzXoqelOSQ3VgfARn
7cVfWnj/ayt8ghUPdiAbutYaFKMzEaMHZgt3f7kjYAo9tKLziC7JRjF14f+nDlIVGBCf5MaESg7V
AfflChrFFf/TkoD2xta5LczTza6Ugk2vvzyWJAmmmxxb3HyOwBonH52NWAmRcxQMrxCzbsCVCTlI
4amBGB62fQvzUloXPNnzXOGrPyc60DdUX6qgaDvEi25l+IKkeRwbe1XidWD+1w31R/K+aUTUPoG/
NJT4cWWoa6Ytq+9g93h1IXSHYUw0MQ84bXJxIP533C8wlt/BnyOUpRnGrP09er59IGi0ZvR9fGyA
kf3HyKjr5d5nkG4jJuU34R7ckKP/d0ujWgxafBFBegsjq79LN+l6Q4R1uPh4gsJjUx7FggBep8i8
ZRYhHBhpAdONORHTIEhT21xMEQL5SkG+RfrDJc8uDIrUp6ncckk/LRJBJChNNoFsox7uiJac/y5n
XW3RH7N4coCG4ECaBmbVQKEFM7EXjqDEqK8MapoWIlMFLr6oI+QPujXbEikP+RWGV1vbA7ggJU6/
itd4AJgB1Av75keR4le7xg4pK+wF3cTZZP5z7JSJMyttAX6o96keCsitcuSCncl0/3fV3o2qwj22
1+mZgmSHT0Qa9TwwR4AxqQNcXtyKhDo2IwN2pg8PWpFF9Gq/Yt7selOb1oKABI/XPRfIZ7PdIYr2
hJ0pQRFI9Mvgnyj5z/ZqK7dG+A6l6xtag/uVz071huhy8IZ+C/xB9bw/P92wwIGL+AVR8xtE1eQe
oKRbBA/8LSN/B615/jqLJXCe7Lb0YJStAH/9yxF5CLTsJaAGccMk28IFMCtCeFr6Rc7uovrC9s/h
5oR/6n0KL3x3boJbeg/yXYWcZf6PakOoTVG8DmoSqJf5NPQaGCNniKtyorKc99Fjy584Z2k8Sb9L
zzZhm6kpPSLMFR2RBdAtoO2e24+eNLMshOCt4fm0W7Q/HQ1nMNhO6G+oAeR7N0U7d1nJqVrPi86O
ob93jAPmlhv2/hxmn7LKvd79hrVdEqc7W6o3BAjU+nYMe+8KuCrhlmqTgWTpX+BIg1mCif62flHF
FBN/UeWCY4r2Kytd0j2U2ISaOCXX6nqzExMkXCpmjWVisqPSulnqMvaUhn7iaQwDQPyXZ/M1j/RT
SbQOck8u7/7U0fdjdooL9A29yJq9nDNaegSCq6+5bfB/f0IJv+Tkj8Rj0ECL76dPCUWC/9VS9Rhb
A69ePlcbErej77IM1pC2p4AD17V8oxqNwsZAYMSjxrX0/gEjBJ9eMCcI25qWBlYJoentebf2sUgl
4W3xfdNNDgkxHnSUb4U83W49kVXI/FPU0RGYD/9LeSMAdj9mO7x1IHtbkXBAu9jRGhY/ZJ/fjRf6
TAa2HMMUgXd/OIUk0quf6J9wbNozMJOSq+mf8bZW3hpz/8MjmzENWDfzleX+ASAQ/+8nZ/zBpmK3
bhVBo7+so8KcG/GC8/hQ1h+M/G5fpYflhzWQSuwq+olHxMvGHy+CXpe9Jz0K4ZWTwgjYG5y7n30k
eQe3jocbKqwmsCgW7Rq/5GIcG4MWxsG6TlhIFFMkHTD6/5tvM/Kew6LkQm0l+Qj5whJbdu74niBr
cs7gQ+btTduuzDjAMn1hNDPCCda5Zblw9qXiNMN7pjro4JIREKtwvMLfvTczSE76Siqy1AzZOvKb
YHfn2GI1MHz2VwfpA2mt3cxa1pbuj5xmamuEWzoXWmlpdazFu1pKMEPIMLzrVTY5ue0vbbqlAH2o
g5IblAIiKip50ZZryZrX+ig3a3sKqC6ZGI17VcX55CsRIZIES3K2CG+LjmlV4c9Ltq9yqMfkH4Up
5EZi4XAEBGjy71vbnhUKsJP9N6MjKKkl655gUJMHBPArReWHI6eyzyInaUkMhmiUAHofq4NAHbOm
Aj7aY0DM24DPfdAZaFffPV6wwg58Lp2UioTr87pQ9aCesmvmkhIy6O0VTjGq9TXv5asPPV1l5D4U
0dTPB/I7lN2j24WpAbNI/xlKoH+RnVNAqmEPbwQtg3COGKR6SR5HeNjth7+av5TkbGsLpEhlMVdL
jx/lkSa5pdQ7CnmwH3gFY8zdtDXiht0ZW9zacbhvJ8UK0MmhIdIfi/jQMK/85Sv17W/iMandY9SE
Tolwf6FkclOE3ysJ40E4XfSco7LBOAdWBeRan3utHTqMOgxDoe6Cd8gOpp6j2hs6VQPjWjgFqEvz
9hLA/M8AYSrZiLGkp7d01I0Y8XaXVn61zRVEcFf5HQA+Lz9eO0jDVaUN9DBiL2n62rqZ6xPclw9I
PZ2jf3kTqT7f5tC23oA5TNvQDhFIDVgGfYs+LVsft9WLtyneQ87gAwhrkqX3AawJ9ZDcbY9wMctz
CKnKI6idXb4i9HYNZQiSCH+Ktlf9TnmTBC0NKg5b12l7N2wcbHQLM/bV4/ODdQxBgMKm5HQs9ovL
Sr7t8cU/fBMw319hwBtZQqaYtQrkKkeR0FbD6dJRPAoaIkLCQQXXu3s25/6BE+nYZ2dhD3xDtOHQ
EjPEJ+7L/W07EFqQDAMcw0d/xUuJ5Qxh7nPp92+R/N2tCO7hUd+1u+5WsjjxLoX5dqG3RkbGo32w
gMBoSNHTwpV7vjtsgaz5Hfo/XGYW6j/sZeiLRy3Z4RI+ZJPzi0TlUf5IiFUgvmPSVZyOnK9e38tl
ML51to9tA1ELoRUsoGid16Rs+sH99OlPPRwKPbIxYMQ/b4rKT1AvHXbyvcP/2F0f4g5dNB/HUsaU
4JLrEOUUJn1/EqljRmPQh7BzLhUrWA8tOMNPBSBlb8+xmcUM033lwv9T/T7AGUt/VLX/xuEzJsI1
Yz/ihpAVNKaLFLA9oiXo0U8YP5ILhaEtLLZ+ClnE0O81qtw202B4RECaufZw95Hkwk8JoLhqHSAh
EtPJEfdJ0EMChu+ex3wDMO4E5uolkoT4t4LDlZh0KatrL+0WGFuUZEMyqtPWyVqvzdOW1bazv/FL
VppHHtFdfsbfWcd/2BGvCEiW4vYrO7vFOo089AVVloFWeG5sYxsdpyTD45J8DN/WkROXit7U9wl1
dJEYMShjxioJXmhw7l8NfcsVwfH0ylAVUpYpbTEPA6b3sqfwBxLWTWvvQiVRSNAftSnPwv/mOvqB
/4J+YIY3p7d1Kmbh5xAXBz2u5l1iNZbjFFnShrvBpdZFktOOfCefdhvgwbzAtHBzTtoXp+hgFsTc
xKy7irEXRkMuKd8rbrCgbYNk3sI8V5NVY9EN6HhR8MOOtPqnJPu5dbUONbrIEr7SsmhvQT22Jh/O
4nOONBtygiJlR5McJmEBL6ijHNnao0CNkwCO9WxpnIVWKw2EsqWNL2Cpes17U5flVV5LhXIQhmO/
WY5FdX+WtsFI22cidV3GUAR76J+h+rI6yBmfpdN/BLOtPYK6/6Hz9Qj9PCnnTMjiMJ14WR1p+Cgz
ASh2cokL+ITA1+66azmQe2GNwwLZkfv7IoBR0/zGiiQA2b1cxCUEP8LXMLgVfC6LXGvhczLoceru
suDjW0ndT+Lly/H/3P1TbMBjXITxdOQ9OwmSO8rR8OzMe0ESstAfQHWiIZAEIt1SsyPcd215gb6B
6URI9URSA0gz/RH2rpUXVNFPfR0RdQCve98VX4OrtNYzWzcuHZTqjn8Ig0/7NSuwfwgx8ighurh7
ZXhwIWiE3ohImXMwafBEQH0v51N9Tt4MX/2O+S5N/YJnOkq7qxBgv67z+X/hbNUvbUcgV843cjqx
QHceCrNdivILFITejFUyAak7CK/BFCsFW9cHygdmw+mHAz1ooW6NcPkCWSzJK7P5Qp2DFGzdo9jA
2Uh/Fct20cyjWEFTIr3CKWdKny12jJs98/Unw0vCLFdRfaxVTk8wsUPBrbJw/AWN2B0n7CtnZKD5
sYN3z0HEoTvyrSRTviT+4kWiVnjTFv9581QaiSj86U5QKBCYiUUGtsHXKqj6Wu0IzfwWonLXQiq+
9vBY9ysasePwaB2wZzxcVRUSo9xuEkUEJUNEulkPSPs+9hN1t3UmDsbaiPnNSOs6asAr3SmMxTOr
sCDSQrkXsk+joMELOOvGXdbyjky90k7HdGkkSq1FTs2JeUyo/tX3ASzpWGfKWYYmnoYNVXwzadg0
N23cAt5eY1d6QMMQmgd5CG58iD/BurtLOxAcMkBF638diib1udJ2veJ7tl8xmg1C9g7g/mnuz7sy
fFHK4NS0uk8geNu4Xuz32yeMj3fydpg2J8Mp0BoSBrG1XBxg3Lz/WXU4lVQYbDAv8z19Ds+Ex0Qi
GIB9XpJZ8rPoedxkdXsua79I4QhyxUsmd3KTyppi2OuJCy7utkvj0UufdBy9xNiDcfk1mwN2B2Om
jf0vi9sTyksF67pe5J//jI0kYMrUGb64GUNEo64U8UBcQ7oQplRwF3zmhQ6Dh4EWf2tTUO2Ehe8W
xaRVTwDUL9qPr+35pozrotDasqvt/8dGzcVMqcTE/ynYgwPdY0re2Ut4RiTPjG0b+QvBQUVrH9DL
zVwZe9Wl1Dbo6PKX0tSWpIIdqzjw1hv6tcDc9h0wApV4C9z7vo3r6iC4bjBXDd8GTr7Bo5MLXiG9
c9z7YARI4CX5MwoKfh2kQr9mMyprpmH5PQMthdEfgkDvB3rDCxNgsRmcQHxryAs0UkxH0R04BbYi
Xaru+K6q7byNgDzUYxAS7N3tkQUIO9xkeUOBIbbhT5ATS8TKsrjYTRAgBO24ZhzEVlYpA2zMPdfH
ht2fUNyVr6AHeUwvmsiUpqrcTu+B5lx2cdBNMJQauaoyo2sIPm0cM1VpczLcHjTa0nv2Ew6kM1BF
iSQ9i3MdSFdi2nK1rxEtiYRv2BqiX1+0i4q8dBOP1zsTH4YFXHGY8P6kMcdYq0QTkRBqOd4WYxXT
WQUgOtAOT+yqxFfdKPk/N7v5KsDxI/GBSah8lzJ9FwN5sZphRODPhAvzeDlSmrz44A9FJqNNSw3Q
Ul297nO1QTfJlY7PN3iA+5+pDAZMkztHxvzsHjqGi68SgTqewXXVTwDAU4MCT5iH91xYc/VAbMZt
j/pUuVc0LU7Mh68QCJdys7qW4+LKjYI+HJFMjvHMyRvoTuM88ecW2OxFPnP4VkuXwt/yODb/5OvM
RFnXhbb0tQy0Llb1Mt0hWAtJEbncnGARD+1XwRYxOvYuDHuLr/pb3wdjWS0YatoEQhTVeRg3CHZg
MUfVxGjfuJ9ObTnCTejtf+uJI9IM6a5r94UvlseJUx7pficyBygotD6D+b/vBXfhtTHmBEj4sCCT
N53L5URhOKOGEArT5IufLwW/pFE7qyODR0u9S+hiEwwmwtXwTHyLuMRSs8BDUQOf/+qcU8jB9nFK
CWDnxPC8upuq/cSaZ3bv9UO4onEIOxg7wllzTOiA+uwXW/LLaD6dMs5BrItItun/M1CxFwr+xmHc
4bj51dkiimi/0ExiVN6XKdqcYvfG8xoDlHGWgnKie7FeX6RRf/e4mru7VYdSE/sUaUBB7HKYcnHO
NJYfvaUrtbGzbyukBgRkm0zbOCeE2cAthfCsuLjAUuqGw/r65QuYl1S7BW+cD8uO3L1DxZ+m/b/3
RmxaiYvoIPVm18dgwqbvRA1zxBaSKtUM8KTDgxv5uc/vG06GClDrNjZ4y4UUA1wMUELNzE8MsAlZ
wzYUbp4XORV2RJbyTXif26I8jiJe5ffdaVnd001ydlkC7NmN0mqMkQqDiZX4gBTgh7Pto/dfJO6K
4X5ejp3EPahGatA5tJJzx5shpfoYgBNALKafGnfsc0WG7Y4U1n7C1A2N5cK1T0yJc+WsdXhyHyGl
sn/rF+NU5bCsomb/EMp7uCJxpWOQpn7a1rkIZ5dsvVSmRG2DymtNvMMto+0/IbTv1ISJschJk2Gs
8JxCP/G2sOyv9FDMwHHGrgOkSRJad68ntPUEzaDZWnPtxHaA+6ItM6L1BA73x6BtG7hHO9fKE3n1
1pF1eqD8QWq8NNrpreZqEjmAehLgY3HVMBELZFSemgbnLJ/2QVVtZkTvNBznfojM88SewbskvdJK
InRtgejm5LIXS72xuqVJQjYphGBe47j5xY8kYa1m3JhswezIvOsrVM1c9lF0utEuG5PxRxnqn9eJ
dZ7+VCJqzXkksE5TZXoLWUJnoq8EhE/37cQzz6foAtoPypDeANSaiJVFV6dzbpTP/HE6Eg1OLcxM
S8teLu5W73Tvz6GCgacff7JWY+xNcAFwZMZ5xvUFtqayN3FHNHpZ8FbH41ZqOpvHbFxX2IQX/s//
Q7cI2cXgblifWZI8kGl1jC5inwMyVY0jiS1Jgj+OwU6UY5GfbCELyOdIyxN17K33khm6pnjDDy43
F8J/3gPk5tbRi4R3JSkCXRABinHyPbM0VMcJ35wqrmUWs60Of5nxFsA7NkyZpCsm51LIVIS1SnKb
TpIHMQGZzzdvxfDeT51I2ocUcFTeZLn0wVFIMygpQUu4nJ3wb+np8AdgeWxvte/qA0BhAQL6FMO8
xwhPuOwUTaflT25rUXNmrbihMi9Jq9ETbEgqqfc7zqP2Vty2/2jOfOMrWvJrxLP1SK8axa4DI8dt
oRjUMwvMrmVvM34SInuHywEeGVrS7RAV1yuePlANlJ0FblUl4bDxDluwAZXXOFl2Q6tW75AAc7NV
8muyG6xiPLMjqU7Cdv2fcBaqib1u/+mR9XWeMkj0L0J01aQ1FGV1cow3/pWyFJfgAPK3smLxTUEi
TiXEx2JbWX6O8Va2bEAST3kbNZsqTRRQ4AV45g9IBZku2YBY4sQP4uku3/RiwB6TxHwSSrfip90o
6ITWJMgGUM/PqOsZG/rh/1Bs43fQLAyL3iPKK+p7tkbJYsZHz3wswLVS9/fp87HRN6IU85AXJBOf
km5b2+LV8rieWN6Prj2puF8xajswd4tx/DwIJBvGcO5/5iRLG04InIfh+QcA9opAfe3LL8e8HtXP
HgBvTz1sVPlLiUNeE+QBdqo/twk6LjLCJqw7mCryEi0++E8RuGQuDXTfl8IYtsLI7xtrtDc+lCns
WSVpJLeGM2VfbNBMPcZe5UiyxpaaPZVBTaPwb3RRYs9iOoKbnC38IoQ5xDfNDfamvbpDEreayuFb
peLsTDiqtpYoxxunilD/pXaPA33IWW+bO759xNl52DaESWeA673byz3aqs8EbYN6xiXrDlFE3TMU
M5b6LrYCu9H4hfFhGPRhIUoUpjEOWp4xRjgQcCrjeI4npzLB5CFTY/1QvXTFRlA/Cy8heUG6zWe7
chM/TKQqFbBmCBoKGlpio3jah2iOzA2ZF1t6OjBEefNW+htJOXzVBq15NQMcNdHvihYRnzK0fq5S
wzpLu6zl2jkdFiQAMqNt8s8XFh5dioE2rUzmPFcpLVd/SbkgPMEmxE8gJek2l6/UMaqrCWMGdU5U
Qei5w+7T30rYbu5d2rFlb2iRxY41bIqF6/BjFJuqM2K7LvoRdWFCKHjQnJb4a7pHfXHvUdwzieOH
L5rKgt1Xh6V3a1/+kAAiTbu2JGhIBsaOMV2HkFmPvCF0bFttYIofZozGAt7HODWPsj6uQLnGjSy+
2pM9d5ITnQx0nzBxd50dPCWAfdXmDpyzuA2TWGH6M57lLWSItzE0B1dMsFoJBIVICqCSltm+aktq
rdT+vHBrxRdgSBosSMviRG1hqxQ/Y9SmjD8MBzBhJl6DEitkHHVvgAq2/+NElMitDH7Sutd0Bfh1
msGUvBzuabhxSJkdiz3rFOr2Xpee5Sgqo3YKHgC1KbLQMWdFGC6O4illTq4V0Oh5aREn/Nc19Xqc
CXlubz1jhghDAgZ1eFWOEaj26QxByQyNP2fs9HmaOJmXkczZeGbdFfSsANP8Yan9cf+Utl9+0GUV
Fx6skxR1IdZyVTSxS22yPbccb2iEbrD4YDB6etKmh9DJpu69PM9xi6AKISNs7tVycuGUp0f8TK9o
jLBceDjeFpWSF8VcjRFwp4ePhBExUVWNcmzxmqRy8CoR1jdOYC4OZ7mp650zretwagqmXtXsVhGq
Io8sLEF9/PGca7fgKELBNttNQpyxzDdidSb7xN9KlVGUf52Ka7LCy/b2zXIlBnY2cONyfjmrpEsS
TgPVkLU3YYulYhsNaFHAk7xnGdReAMScuFSgcGQHANXDWHEOo8UkoecqxfaO8L5pT3SfMdFzyO/X
ZRlS6Rr9VPLTo9L8uZdOnmIedkcOV5ui0cbaRAKqdQXMS/hBlTzDb4fHVFD1J5THTVeQErNS8ZhP
QvhieRCpaqmYEWCgyj27fxBhvLlpOzzF8Yf0EOfMHzdeZ/5CA/ejvr2NlxczwtYKoK0fTowYywVO
KqF8i5V1WBTGWD5pmA/SHCb9BJHmnskLjC2Nx2jvy97G5J/Jc26X/S6eK2g8JCfmLAVwX9djqb3X
TBCfcdFBSU8Ugn2wXxudXDA+7N/VNLy39ClafGVMYsjRKWp71H/3ba52vIw6XwFYf7BtzRM0mmlT
hkXA5c4b7seyYRZAAmVu4aPUpDrO/z6P8oMfzENcrcxbKcoI9OcagodqAKoFigX2OlaMSfFmKvhJ
qBC5V+prVaaPhkozhQIHA69huOhj45WW0ax6FoPkMtQYh7I9DrGQsMgbAwgGIcp8vc7WVW2TI3xO
v4c2+B8+SqI2N+uhBUZtH2rbZsZvhR2tMK/FR4MM5LCSlDF3Ase+WcCELediWAtdZtorFyZzrDWS
xre+B9f20Ab1+oY0SxlUAtxyI1o9cdwJWYGeALi0Q72DB25CDAPujm70OFfTU+41cqjiegGW7DVi
cnV1+XAPeEwpffCpgDHFuz7Vqk9A90xqzKEB+/RjcG23GBHO1QiSwP/qvtws/kOtZUN3AWA57YUm
5DqV2nz064mZgo1O9uhnXECakqAIi1lZ0CzWvB8GCOWygZt2JodRTgieUj+V+YbLThz8wBO73xBc
GiHwctaodxcWamMwBvbmeD4/SllPNK5Y5FCNP0xlYZxwwO5nhqnYlju+rkXzB0qUNJP2GrhppHE8
vyFX4YfRqvERufCOWmERKYPCF7d8WzU4LUnZi6pteLrIlbbomyfGzsbu4m+e3sumUyihnw7R9eOA
mcDNrvR9t1oNO3OkPlzNThYv2XnfaZp3DbciAqJj7xP2Yck6wuHySHy5xAATVkcCvscTi9Qe96Kd
FVyraTLah6+hC6309CMuBW361qxMEiCftVN2Qi5EsXrO4KWIIANPHAggJcO1MMMXGwiwtJr0LTVl
cKJzTCVzywruRaFpuucnW47Hmm1q/SNZoPAwdvLCesUpv8XaAnPQBXqsOZbiIhqVXyKq2Wa1J2E9
WbCJvj8mSR+TI3NrL+v91qzsT5kl8q9ePJbTSc2PI8GPk+pmDu7dD94xeSBJGSGdURPgKbQ+HnC1
Dng+cmdSJDeHaOxIaStoR9l6XqzxzMNcc6hmV0joUMpNsZb0h6c00QLc/JmPSLgbgAFHUErmUzo0
OSKrYnFuGYN4BqHoLNSqghj1Cna4eUb4ji1K7o3xgnsfvIDuYm8+dsG4/WyXpz5RVAhnAAH3Sxep
423TvFlhZ7AJ1APsEA1v2NolOnbIQudYCRWXgAIowj0TuUReJ3JjkNCDdv2MI0mAPEq0noAs6py3
R+6quhdrFNwQge2P9XxZ2PmiGrqhYNOCU99YAL26KqJ8eG6ZiD70yVJGaas1llr0wtFs/L+19wVg
spb3ZVWnMBbvXE4ZMiK6RkOvTq3IUS5bU+nECxiuEsy/8ou5x6SP/4wN/azQrmdqpqGIPm7NVjZc
uFBMg4P2IxH8DBx0+E3RlKgmcz+GAzgmUPqFeAEghrgif6jyDYFlgnKyOphHrqm6d3OAWPHILxXf
X/IyIX+rtqQii8cqxLgbIGKSId9VGFwvRsFmXH3W3gyLpAcgrga65E9W6M0HFymYH7VA22F/d7Au
28KdGou0D0/x8W7GpmUnZPtY/BVTVCISIApoqaUk6xYmIduuOMg+8ekqeEEqrulGgs5jUKhdkRIe
7eSBN9ooj/8nwgncOqPzFdPQc3F+kaQnh9pCo2yy1GF/4uUf/Uc61Ck1nlXJEmiRp1siuU63cbC0
9uG7cXrDdZfjYJhqdXfwnbMP640s6HlvjlQcwDUR03BiMgm/H9QPOoFuEvnrO6bwDMahUiJUaIuS
HtWVRo0q+NU981ich9eo9d2bU41eczXke8NXXpbZ2Z9zwEzs9k+z8Ro7iMlWAvJG4UN06aQUDmmK
8NgICn5JT1V/ldxthxJhnDLkla2AfYExK7d/MN3Gi0DQ01xqYLLwW4Po+kY4HN4utCsdalDXQ2dV
V8BrBcx9zP9mQ9SnmuL/8oz1xOwiM1ejY/cjk19sTgnRKcgLJWq+qqpeNxF1uHlPjZrd+DVq27AZ
xQU0zQZ53eiM8LOIfnXDwgo2Rt2r/1dbuSf2r1Z1kTP5zYm5CGPd8vMmr4LH1iPknilGgE/nAVNb
Z03SaJwJK3TgzQcDuEp2fQXA/dl1ZeOOpgf0OroxM5gppXeh7SJRgnnWVUl2WZwNMkphv2XNEGzh
hNix4LLLI4qQGbgC6WIMmB+5HyzxYi1Vk1kssZIv76a4JV6VdsP5HzRSmWYXyo7ZmoaL6jT1NSuZ
+jMrkx6aL4JMVdFHrqakx8AlxmjGOwDanuv5o2U1cw+Tn4XLa006VZYv8VjSVfQIMIh0GaOVo+bq
4fzlaZvmmoGY/410K8C/dzgXHlXcvzqEMn3/PyGeuxxlQLMQR6rDqxZ5sZdDfan5JA2dXoEWnPIu
CGoaHlji3YVCiEScAtHh3a4a9L7QSWBddxE6RnPd+WLMVRQeqTas84BTwm2C+BBC9m7xGRvfkktk
BOSvFtFgBM/JV1ii1xWqgsxSqOzVOlfLFbnXYaSWuxRcHCqCPq7rar2FRY88lpyNMUB6ZdigMeQd
itv56fKYRIhDeisXc9QgqaLEjjGO1JZVvXrYj/H709CTshw/NWF4oTSi0foC08rwQYusVr5Ut7p5
dY/CKHZwQSB6H8x186B/2plWdSZaAPOaVlQ3vMZDJefvN/PyWKtCL1PzYMcW4ODE0SH5RE1bN7PK
1DfNrLSwHqNtGxXk/lCLcr6JiCV9f2nx2b79VWvtPpNz+tSkHTB2uVXgwd1MtxQUCxkU1bKEYQEl
5LISGBTwIi9NsK/YvXk4QnIIGbcrc87gUaQHxUcY2G9TYClrV1VCqHulc27aD7VreaTOXgTq1MT+
fQSyxfzPG/kLM1JRR1XMjOSioUCSU6pZukeCRKCgSnA5PDdqEMm3m+BscWcWOSeyH/WHLk2cHHSk
QTR+xwvMqKPTh6/syLlAi9n4QBPUD4pYi5Lj+6WUKifay3LMtH1eYC5Zw4JeDBVvA64C0FQ789IH
CnC15yFFD44HM9fsbl7kgjF0xlmbxcWqyXZO8RQNWwySXn7rdGsN2Ft+PnTz1zmUezpaf/gGI5OJ
DKtT/b+YYrSK4KwFZIqDH4hw+78cwqr38x9OekD2sc9OIQnWTiScOEFqa9NYfAJFZRaumwik1Zqg
HRDgXXz5ieHIYPYiO840PKdt1r+CLeCISE29mD8+1hKwC44STLabyRxa8xdeKX7y8e/XMcdrtehf
Ka7CHQu5NI3KOrcek9ninzck41IS0/jZPHUu+GZmyH0tRcoVjcIerTXrFvBFp+1GsFPIGxrqXSfK
GORITtq8FGEcc/bseTLVk8VejoKyB5PNQzatrYvutaH4yBpaXNpOmRuXxdI9nL1lyc1ypqUu4/V6
cxPj1J7RTsUKah7yxIVYo5SKNTktQTN6OZgfhrIVFz/ybo60redTUcCVObPqrXnWVwDyULgRVqHo
3WjyK1dJYl1sinoNMeeSeBnSUgzcd4mPZp8tUaZWdYcZv8ks8sJcYmFVtM6gYai6c8OrZZ1tb+KY
SdgaAETujHcLhlSfUafBRdAkKbHFDKv7px5grkf+19b5IoHZhJ2jIE1GmCSL5Sd9unI8xdG/AQ2I
gQiYnn5G+4Bmy1iyISlpV+lLanzsmTvdGLqcy4/4nVVsJsIqXq1yOIhpBkJcEjQyxO+GSpx7jZ+x
U5G3wqiFK4nbUeYlEFNoPoVbjeHtZx310ZiIA4Y3quUeX6uSOT+8cGg6IB2yWFTBkj8+px8WhI7v
sl323jARWLYnkUjhuPzV6HSJZ07TfWR1zIiKd723G1kfy7P2JO8OibZ5P4IQhlG7imRsfQAlYgUO
kAqbMvA/SZGA2C4w8aa72Yrj1wQwKiWZ2cY4T9OOX85WgZwkrpxBqVgpzmRZz6ZNYB4b6QYDctMA
8JwZLfF75ACJn2b71Es+dWn+EYVweZwp1L1whIHb25LhmypuLbyQHiJAnCYXUXEMAoiu7Xyr8doM
nwJi1Dcel4H31Lsv1YOeWBWbI5PH+YT3lJ3Cj7vaiirOmszVBeWaxmVoOugU6o0sKxApdkAm7ZkB
5wIPGbDmU+wn8fKox0ANWClqo3lYlZDx5Fcj8Hhnf2ommZv5yQwXfmpt8xGlk9sVl2+dY+ChkqR7
uFhtD/gmFUcsoxDW0Xc+rXsPh/j4795W9s+fIg6nEwOnULZKyz9/8rWLtbCKM8GvYkmpjNMTzZmd
qQMtLGO8G7Bmay+f0/QtipcLZTHMH/tqFn4CEYFAdB5jYDgyOtRhCy4z+Lv4He6S+bNjyzoEuWGH
f2vuOs7llSh8plZumVljAf1L5CsauWRaQm6bMSuU7VeCwxMEBerqfDIPUytmISTMyNSPYh/iJuz1
yRqxEOGIyLRXyh2xXeYrKf0RyL+TI7xNdwH69Ih1eFYp1a6+JBNqsdAI3PTBbZfD1gTeVD5fpwTn
fszl5BAK1/HveTsV/UD0EA4kf/lCSDOtnW4+cW7nJJGu0iTpkQ6f6bGSe3cI3mYiZOpfv1bnJZt6
g1W4GA5IXtcV+0Uh4ajtzc8lUUEBPIeCF31u68BNvOwQfBErfJLhejqzUeLgChthFEbeYhAYmOmf
audgr3ALpfYwvyTnfhxcQDlD/2z8Fy3p6OnNQIXcfhWd580LGFHLdKs5cVjQ7OMUKSk4zbHdglSW
yJn30XAH8PvrxtifTDba8jwx6Oey9NLyUKtex6/3L2zD9jhFMuMUQqmnIppLJIlQQ3qVed+uIStT
93m0F0LWBPyAQTzmL+5P9ok6J39pRhQyUJi3oIF3STTyVnwvq4wc8T4HhNCMxTJSW5yN37JQUQV7
7Ex5uMEmqDzXf22aWHQXkdLdda5GMYtFp0y4PUEZl1wmvFIAuRpQLJnyjnQ2Qz6m7KPSXGiab+8H
oeEu/8GFo7prWc+cC5K+nS6xe16L30+Dv9AtdNKBCf0cvglgm3Ej1PZx3K4jIOzebdDmfvZqYZvO
wq03bq2xUpmqHWEtG/uqmAngxNP3LHYbifjzkAgaZpMyKwl68AhXWlkbdeHRG7vV93XtYtlPOqDD
hpWdIxCYPtg41VEKeu0Yiygr6THMzf0lDIvc7z6OGwmVXP0biFOfqEOXS45iiFNjlpZ4IuzapPq3
c4wxcWqTiEykjzgwAAnYpRX5y6b5rhepjH3Vc8NAmsHva7pUIcvNIwqP0IwFM98Gk9HYDEyu2H1u
1hcdP4Rpy59/pvGZytYIHEurtroyvQfvYAtFr/Xy2IuXY4rxtcaDfSH4OM4ydZ1oYRuOG8vOlt50
0SLd92wk4aJBt+g8Rxn+MvCDecI6PYq7K+yBMebRNXhsVvjEdK6mR0AXQ3XWbmtLja6ZZfAuejk8
R/asUtSKZ0KCtXZHXYS7kNfUwtA1VGIqxtvlTtwuZ4/Qnq0eVbvEZMi4CL8NQ2i+iVFGziSl/iuq
JUKrMYe7BbyNJUiQ9OU1+opR4+hKjKdcPsO0KKu3Z+ZoXOHEXjnWzbpAW9DhMw3BvQjWifYO1QKX
B00K4fO/dqnUw0V22IWpAsgCXN+mLkIxNPszdzdohPkuqljM/6T/Fo+F5rS/YrJ1hIN9Wa8xUFYC
G+HJ93EJsvbsxRIy6g6AJwTHJabrs8JIycstDLr/vDcd1RWt+XOudzWiiENWRSnXWP6BQFqG82br
gzBh0q90RJMacPtt5F46qlXILJBHpdIdfiPkA7O0o7ZjbMYYuSFamly3gn9XviJqbK0mjQZtU6y/
6RH1793Uieye8s8cT4TlicUgbQdYRqy2d/04KFvL+XSKhU5hDQwKY3cZxQLQXaQT3EeULTkCOfxG
yFYeiUdxg148j4v+FdTrwM5fQXfXyFocwwtpjc/Mx651lBX4sOJFZIGdb2qLrtlvufFYssiKyybk
A10YIB4D7YqP5dfKFM1hcFVQGfolydQmRWTTQTOWmTq6pD40mZd7tkhTagl6rO+yT1wyfjrwF0cz
OfCxNy3GUxhFbD+B0oGaOcseqBFXJp4TfCDAyHm1gsusiWm/u30J7+yL47hPpRUZho4wVx5g4pkr
E6woop+ZGGclLchGo7x9BUeer1Lrcph/+dTgrQWU5d8GX1yjiSdttmAOXOQ52+L477sAXH0d8suc
IKN0wvZevLbD8/0As0U5sAZfv+HctDbeBN2htiaLWf2mb/TndpZW1We/dv8gj/wRJzP41t2RcCOx
8n1BQItkSiYh8WIrzdWjwzwE2Gp3ondD9fPVKXxlL+kgDnTEAoFNX2M9EJgOgfp8PRp9iyDvLhr1
wguLzKVnW0LYkmJ7EjCH2V3w3GWDYxB370skUsk1Wyga56uCWTpQuLmqY8TKiuKOeNPcKeG5uO0P
IBxVSIbZdcL0taHepzPyxxPrCK8YqTqNMLwEYkwugir6MYrvLqwJ36NCKsJAuRL/hV9kw5BZ4tNm
u2kAwNIbCApjxBAgH84JdvKG49Iqwg4cJKNed8/56YN+DPM551Uk9jO+cdTHRa1XG6iTum5QVE0t
UPTsrk8UTVQtIk9Bz6VBF2fkHh3dc3rQX/13BuSN04FZ31pXxekGYc0Qk6+HA210h2L9oNvJ7nEF
gT17pN/tddbdZL5Y81KY93YLVj+AwLUqj1dxgmOrDt8FPTNfyHyShpfzr2WCVSuOVlSsYU0ajMsD
m7snszC54Xw6iMRakBlwytq3YiBla3WYnqOKbFZTNGsfr+JSvSH0kDSzbFsehnsFdzuq21dmor0l
eCOzjFG3Zek4KYat19CK+IYS9cGdlqZ7QmllONg5cwKklBsqTDtSE3MFusfyGS0Jm7vr3UibxnHB
C+f3uVMbY1jWGdcZG+ZD0Rwtt0xOoPyoHn3yPpk/LfWvNLofuzG4VZ/ubWTOQWE4DswC8A049pAb
/v6xuCkjteh6QL3LCMJbe3a9omQOeuxMTe2N1/MajMC72SI2jGVAy6Qp45Dg61hU4XoEevNj+BuC
Nr5/U5wsVpw5MeQ1BB9th86eAEXkqAOae7v0XTqr+v0Yr4Sz7+BTZi3rspEjXNzIFmvaJFTO1FL1
2Cck1RVDiPd+O/NY6KXKJ+mccvY035qZ9tJrD2Ih82oLsAmClxT4IW+CLyVIyg0NfqmPcxlaLhxP
2m9AcqaE8yzFVxUhKKi14ZpS6q0+xsrtN9nuVzinrXcxfAn7s4ZlspcuT+ol1ufWyNubsH7fkExu
67wFKIJ/2ZAPSX4yDlU9+LE0ObmiZK04f+ec+7QlrRSg5SFKMgR3gyPKvBtquliDEiJATWAPnkh0
doWIAvQ1RUhx2ltv5Wu2cZJ715SR3TU5ijnPReGhyLnjEgiIHV3VAABkyP08IBBPnbPrz5qGt3b4
Irv+uYbZ05OW/7zYBfBsh24286MciPnW/TADBQz7H1daPjElattKjbvUKcRvnMihXRKXkc+cxXof
b9mDksduuYCrxWuf4HXnxG9/gUhmdiFzZmnmKNx857Rek+h0jebMNAd+AlNyay56hFbocaZ3rSaj
K3GyDmJSaqCKzI/lVlPTzV3bTYFJe4+4AqHMfuOCvfzOWEc38oCsarB6Ze6mhp1epqA/iswhXj87
uu88gZQw8i+f7viB8hQqWazDTeO9h0+7WQ8KR00U0vpb/QiAt/IQdqDQVxOZNv/zBYg3gmkC9rT5
xqPe9NNmkL2uUfu+MrBQlJSbgCzCC46X9tr/gfWuvaRZd5wAYrOxj3kbIy5ykGkrg+/kThII/fzb
oK7SRK77tUuLrM2Q0G1G0ZkoLIJ7/BxK3OCfNnegpkTF7FrAUyNvd/IfLslFiEjaZhOizDX17Fz5
5pW5OtRjJTDuMNKXqTxWtj2Kk/3oh3cVDTqYuNb7BwotcY777Tt0UXzyzQu18eQ6VmKnhWQRuNdd
K0v7XnsoYBJNVlEdW8tmjiSFjGi2xbwBjVNE3mgWrZiiC1MSkJ7Sm4AEIFLZv/KCUr03+uZuKiUS
eNsDA98be04/k3mhv1fjDiFSRbUqutjfUuocXB9rpjcNvW1eQViXYDviiiLMHFPGFbZot6E8LcHt
0Equ2fEBE4th/GycO1HQkbwH4teOsubRnFQ5tqCW+A/Bab+gbEisL9adFKuAhHQ5L8AUsdyrT/Zg
Vsjfdhg7JhKaSwR08BTjP5i2cR1bpqCs1BCDPGIJgjZJVgtBMM6tp4kPEO3IfXtjrxgWbOnSno/J
qPPRabY4S48ZGnYnlKVzJjB7vq64+x6Izfaw9Ac1129J8W3bPMf/+oIoxsTjPgybUAmK6n55uwAJ
RBcZJ/9+b2VUwhcbqnltBXvYwuuhYsnM8XyAzluFv/Gm9BXcveRK4/ALLXehCXtJ5X6/wPcBoZjr
PyCryRpC4keEp/jfMNqwYZK1PTpXr806n5cW92T3J00lH0eNKi+LJzd0G9AkifKYjog+F+dIeDxz
dAiMVCcv5inROOXq/AHMaWGW/1gPj6H4kzVYPsd6b9IhCG3wy9ha7s42O5dQWJaAqHDZG+aeJ2xZ
xvQtXZvYWk0j/oSoLlgbEKVsy/plqN3znvz9vsPa2KtgkKgF8aL1IeGYQATGdXGSYlldJZUTL0R6
sm/ui41aBIabKsmsg2/B/1JtcumY+tfgBYSgTUhjG8ZtyOYb6DbPjmXWO4kLukFWkwIf1I9jHqH7
TxgmKCWOQtz0AP/ZXeE57GQAuTZ2/dvqMzimfiMOduypJawvx13Ne694AfWGuthcvPpMri2f22AV
JR38ndGZx7rjnS6IDVc8Zlu+StNQmnDvGOrpR3cLS/Q/h74bMuUyWTmVO8T/kBgTSyvfDuNX8yPw
rvyJnsLHH4RRZ9JXgDYKLmJeivo9F1sY1P2ZKaH6EAb8PuWZxLpNV+1B3hb8yXASubTAqJperc6A
y/pn/1yYAGac8R3huTIu+j7InrNgdfotZ/xvflSzevQ8cEQx7uD/yrK+ImbrCjs4aZUZo1XdN83Q
aejDRkNP2+3xz6s5nE0X4tWyzA54ceriSuYyz3z8hB0KH6YZ9nTPMX7ndOcJwGeG+q76xPvwWV1L
laJ1vwi/Q0fweTcy42IbRmyudNV8F7BpJe6KJpqZhk8oYi16MvyVofumcF1HkIwvc6l0NFmmrVGG
yB+ZzCaLi7/0vjJBsLOOmJ0xAiwCgyfTo+Z2+LitJTwz2jZn/NtOky3i8u84rDenqHtcaaR6r/H/
wRPFfFzI0UajniQESBbF8kMAqSwP97GT2J8xRNBqYZ46CiDFxAhsO//7PFsYwCFnI6KJFLt16KjT
IbK7jDTqRdAWWp3K+0dkC5Khluc7iYpdJxkM1MbyrqkAfUohhjVeHfReogoyGorCtm93i2y4e2wD
ki6gjmw832q6TJ3NGH1ukjFs0CQv78Idg+gajXl9jo+AWc6I1SnxSAYRL7Aie4Yo8tp11IYyxik+
BRNeI3qvfTpU+oi6XqqnCVhgvVqHFgwUnq+yR7huPtqWr8PTd1LB/zQxFZa7ConsBsnhd3F7p48v
to/DGfyU4jmzpM0zufu7/aP3szv3PvQM4Vb85igQzPiDmjryz1+xl6v/Kba7B/gRvd2pwuyHtUty
RU8XU0qaKt+PWa9iE/8cXsBDjxWc1dbit4FumfXoTsit67eV5UQ35Fc+mCmndo/NQOFf2euv1erD
AHh8RA6xe8R3BV8I9cbMA9fvoZ9awHGh2oqj+4nuMwUJH692szD8ehZjSIerkYR5I2phll92ziZ+
dCY82un1RnIy94nTai7r7TY9PrHUx62wigDcxJUjNbMIrC1NhLvnn3BPi+4dRymB2W21JFfhuKEd
j0cLyn9LBgzvl5++lhZbs7FTFxQfspktdBaMP9m35aaB1+OODvULk+huUcdkQDrnNYfmi4mGeiEu
I7cr5DasyxQcCa2UilqCaEGULrMoOvqwwdIQmYpu/349GP3R3ccVkhlvJy0Zrn38uk3wc7ZyEbPn
OKKX5mGKY1yVbj/RapiexTLgV+wKI+fow4NQtuqCahDrz/y62UJYQQNzUYoK9zn2ggur3N1LjjU7
SHIdJaZE7oEpWc2priK+MFfAK6zYdf8URH9CYNghNS/jMhnVxxqn7pbimFV04FKTLu0j7aSdE94N
NJSnRW98P8uPBMU4vlboXLv0NcG6+qVC0nGZEHl7LYu30mDEne6Bc19hxNCtZnjDwAlLCmyf9ODt
dnFZvbtpPMnioYyFUcDar8fqTapjiQ4gX/VdJOcDtOumS6LoqWdSWXA2caQ5LGUGi6U5e9N+qJIX
kDdtNawI51OGjSMEGML5J3W8HY/q3zZtsTxWpnI/giPM1YC9nLph7/pFDOtt/YB8ymjz7NIrrfAY
8tjTnukYe8kI4gyU4qW9gT104qGIfUaH9S2hgrwWXdbzgDr+zOrNy584Gy32Hnt46vZ/IXt8lHSX
MT+G1Fb6W0NMYE7Nj9HHlZCMtSM4njsdBOYK2JymjI66aQspc0HDu9klyYcXwLES7ztTRYxKxz+Q
aqIEL4SVzuPMCTxNqKdIwAp/6x+tpsqKJFS8CExAMY8INky7TJD2x1EKkm442UBsBlJfyjSfdBTk
7ivw43m+sJrTaA51MduMZ4n0ICWxvXd58uhnJfmGbWMdEEXrj4Wq7ONYZYrcnH0IeCpc61yTaUTO
1P2D2uAtqiZ+APJXjMthHwEb+r9GSNcsMr3UW7CS7QVAZNxBm8sq/7DFIaibap63X0VBX0tnLQ4m
heREFP6lvaozCveGjyBzI4Yh7nK3NT+JqvrXDhXCpRN3L9PR+tz/tXYa7EWuQmtMkZWRpcoYKt4k
AcrDXxKZWx+LMKl20jyMT4j3aqFsc0wthpo4YrPH5XoApZyy8O3+47vTlXVMjO5Gf3pvURUgLPLb
3sZPTtmyp3yprs86WGvv+M58vRQwdFpKZelpx+J00KkC3EIt4Q9aU4usbJxoqkNuaSCpLMyhIvm7
IZQbWlH4bb1UZVOul5DxZCt0Y3LRBbuLOXTucK9TbdZHW3H6t3z/7thpw2vkSgqr7ESQZQITJZlY
KB3rrJ8ZXa42KfPgDHef15p8LwSVY518ZpK+J3+vnStfFQb0wxLiLHXikkfjv/FAE47KUjkidI6D
76REcUjVMWmhyRIq6IbPIIebgNY64wJ15sQhwWkSusjrMylX05aARYPvFrNHvQmDrRB2GuN35yzo
7aHSkHgNbhYmv5eLbCr++YmZ299Qkpnjl04ALbXgLhWxsqCUTakigqWfJ+Kjz6zeNrkmMJLMHlO8
hCxOLj++6KeIDRbDCPtLCZzBHgXrpoJ29j2SGaDBQqcw7rkc1BVYBPvmxZgzlr2tI+FTF2+nLG91
y/nMj7FOSQt9hO1q6uMtbF6zjyUSfAYu5TbqEpQQN1RsCXL0OMbeQxJgZMukmgasF6v6cnbmNyxX
F8ygOmdj+jlCF+PLbzA9JtlJPRA4xVvdw44+asRQx4CCA+cc0CC9V7nYRkvTHnS+Qof835UL4fie
37lD+q8m44EDpTNoHTj1kvuQ64rFePwpSqSQjpgX1L6mmOMlmIkw8b5hale34IRx3PMsnBc2m0DJ
bRZcM4ZeTZ5znyXiqX9MpaVHTT1GGG9KN/TDvqVYc/okXEpj9MsVC94Xya7Q/qijuVuqPr0Kt9Fd
svLyMWBn4anOO2uyMYf+4Ft+kRPx6AoJSmreDPh7MVfrGrEij2WWfh1A9cm9bC2cF22Bb/YtwhS2
dWIzuFjQmaaYV+go48+jJ6QXMFrLpZtANw6R5hT1+OzTI/jI65Q6yIzfJwgVMKiZ3RbligKNfvye
ZcEidumH2Veu1a9SgwiWXskAyl2J4Db1N2lD3uUO7yIWQZ3bEVbHmOTWifqF3ZTSnbAKn5XJ/zS3
Ma863SmRTE1wHDbpMjBiamrUzNGO8ZIycX7pzFijd9zPtvqZOxHagtPhVjFD5B3zvJUrolmhneFD
siwECABM/Ptx2nA0wh0EKtIgo0BtvPBnGbjhOu8yPHXDNU+9MiMusyJBfICFuh4qNGeQfZGFksbw
LLgxd6MloZLYlcSX32e0Ha+ZbCrtF5sH76q/1AlA/ZHukUk+T0Q/sMu2pE9cmkt9m7gbknRqLRGC
6O6FSUfzlMk2yE73FEolexUbUt9QlKiZ8r5PyXLyRIYdp1M0oXyXq1GWMpWHcNELz3pmwuGtUOSq
uH6eaOxLz3+dLJm/g3pk1deXQaFj6ALVCo149yZKS2UmcYSYM5wyIwum64lkA2piYtkvRKYbcppK
oU/YM3lmYFngMIkSlP/mY3vx5mirr2Niu8ALw2OLV2bQ2TdDHtkGOsIQTsHS2N2DlbjvsGLlxOzD
pXZ7JkdKsinpQLEkY3FirtTMIN+QqG9s7IS/JCFwQklsPgpfDiyjyAPluz2OwdJva+L07Zy1y2b6
upxk1dcC5sNZA+oAVvN2oV8Pr9rYF+YmsMJ/01LpJnxQKTxlTQXIX+irju04Pc/DhhTOpAvT9HZF
Npj5DeWK5rEF+wfhVe1h/5e0edaJlmc1aZala8B79BFPI1Pl8ep43RX/yire7U+F4CQ/+eDxc/YV
COO83KxDFoeK1L5Y7a6aIQnc1z2BaN5vvAhkDkLrfxxWxjePHYNE0O+17/reywsaBai42e/ZGcWE
gasyHVahi/W83mMOGvic1wCi+ObdyXr40WdYcuvuyu/gNoT0aJFxu5S5h5etpEAPlUbxrb4x5eyx
GAJmY7XiNvMf1da1GNXupRLGLtAb3NONK22RvEptvLeBk548MoaFRbfQGBKzDIEDSGvQBT8N9AM2
rlgUoaVC01k25cQKcksSHlUCzhiBDhW9lk0oQYrsYjmSsZ8CngqO2ysPt77nvl74Y2/qXuV1NCOK
SwK9jQ1YzISDbEWwKFJBgWvBH5+dAdjpkekytEaLt0G3XfGBSzOptRBwQYZ1KlcvzPwFziF3jVkh
M3VV6ki3dm0w/rwAglH4mJNllUOpSCZUoJqVIWL2GVijVLFhDe0/ubrsG8wvsfGg9Zi1limHAhJ7
LP8v5TGDexlSEZcoTbe4I2QOJ6dcafmaltf5PDabFS5bQOsRcEh943SXE3uvc7z5rnGRlryGp52l
cqkUtt7Km/MbmEGN0Pm9WfHhomspzMvP453YpRaoX32C5whU3hakLAlNk9g559oy6Yx7rPFPrhix
7daJhmR+QTl0/lWZOqdxXwuswtmfthBoQUrYaDx8NeADDb+IHS18b8PdW2CU+ftTtGyacNPmf/EI
bA/9TKa9s5duNTl5vkTduyAnVLwutd1Edyqes3FAPhLlI5QyVBkrOIpyueUTnQv0mLWjYsQ8PPl/
iyXP46kXagj9WApuuR+Y5wX2+7OBkuKY1S9TUZNFi99FqLB4BytefxZtaNbY7SS1+5XsU81CckZU
nLGS2U2qqab/LL50lKLHEr3+1oKLc4X4D4v7VvGH2/v/QkamzF+5K3B3KoNsEmyywFxeel2LgdFN
mGskT7vEIT03Gfp7Tx7iS0BOw6A/f7YO3W8Jctpy6Z4RJ3DG3imAeRdaaESYiVCzPjp5j+ak9T1K
erf4ktLDbRNIqPN3Gn/tzWxGZtSOyuMcnFbNj1kmQ7lxXi9AEe7LCesE61a7rwgCppyWlEe5seIH
A5nXCwyAzPDDsojP5HY9tKf+VsVhN4N/inpLTuKeWCaab9obCH+XHG48MbiqYC345gs+wzcxnQO/
Do/NDH0ID5VktxWQVkq/qMckXVSH3eMV3WuZCh0UZ+PfZ5Yc6QAIpUTvTvLysR2j+NtMKrAxZdWC
GsYFpKDgVP7cPsUg+30SZQakJMmiez3kLFlIMduaokeFy+oeNpJpoNhIWHCSCOdJ5aSj8pMuQM8W
R5MFau7kvDzdThFLV0sQ+VmP2EmzVzDC1vMk2htua+5Q9azhn75JWvSwG9BJeEMGM9jiRNyBIo4J
Vt4YpkhqMHqwjt5gfv6MTJl3ZYWvRIHa5OBT+H80d9dC0uLLtoQ/K70ktrLduijA2T8Ly0z6+HOE
NDlmV9p/4QZlzVLftL+KuLwsRTcUjsZaX+kAKm9FNLlkCzSsRTrBj5Hw8dV6w1X0uTrtQWEtMENj
3o9MPEXsuBhydm0vMPEFap8VZqUkxmDLS6AB80lF9YuerTm205rhIhRZ1rc5ltjEz0m2LDXC6QH3
LF+8+yGHtofqvISSJ3e92jX0/aOIMgBMJM83cHYuamqC+QTy4LkI+3zjGqYUQ2vLm8EDxaZ/5x1z
yr0ZA9JnEK9Zz0OxkT0o4zh0ZRWOVtWwlmWPqKBl9xBQ7xNo8ySzxOJMmR3r6w1BY1Nofy8M/oEx
IpkBcFSCiercgUuR9/bGnM0GN4SoDrwzcEFXI6vBCwt6L2hhPZV6gwSDw03SnligPGSAMLzu/Lu4
qDrq6U2JPCk6rkFjNV6XrhPNWr22fnWS6Qtsm+HlLg9W8/ipNffvUGfQS+Di4IM7ZHyh6nD0UVYq
GlP1D4ZjJYr8mtw5/3vaNk2oEjRqXBMBA2xCCZQbl9hyozoEx0wYO5Ng/5JJqDpS/IyLM3LGkYHH
P3u7/qpvgInezJu4W29w7L/43oOScggxIc/s5oXDokY1ZWoR29KL7VOaYgF8w58FgoAAwg94gn9S
GWEkKM3Xo4tNU1QwUhqZzAAqQqzRNUU5CKpVzMYtzgACXAHA4fwg4e+o9XfdVN4AtAHBq8csJBmP
PkbUebi4qFjOYMvvC0Ykvm638DbjMm1EsKLO+5IYXM/1UcTwn5YZ/sIji65RlVVrsQm14/sgEU9C
VWRY3ZlNVkBNGZFGWwPmqZQknx1WO/wBBrkE/lbDuZ8PHp4hXbMNSPtkQu5hqs47MTO2ciwi+0j8
xDSkPi1KFgpqm0cup65UAczpdPcnYfvDEiJ9u0TeXrVXxZQ7A2VqF6eB84UiaPuATPp39D0i3fRo
tstRwGDD4z40uPMm80AmRR1n27yj2m75KpkHNldsWqEr9wGFboc0NCC073wESTjlOf1q2E2NxRL1
Gs033Yl3EfXoz6fbe2kvCjUy5gWCdyu/xXLfMgFfYtDeYnisYgPMQZ94m3ne/drb2IcYSlP9z0vV
ih9dZPv4lp6OjUpLgO//LO8D6oKlwfelUJXqQu7HtEIChtJ3p6s9hcepKBIgkjfcxYeS5d/gkDt8
k7jQQO3zFWnKWZWn+2TStAW/22dwUtJTxo7no+viapu4JWgi6lNwKNfavHcpPIsJDtzdV9LEfsIT
x0Bxeuj6dK5V+3vdOkt3HQg5lrd+/5AhlmPcMmljGnK7GWDwmj4cu/bsfkVBWA93JoJxiSLLoKzf
eAysw23xzpmmJ8nhxog3GpJFTtKYGHXCbDpQtzwaI3ZknMNLUifcQ7TFY2YOIPH+R5m3HH+9yYWh
rNSqEEZ1uPQ9hRR4ugfN+Hz+mgRQArQ35sQVZSeuhX80kspacwb9SsTPK4XsA68mA7AKonAT3uxT
B8HVEquyW5R0vtVhHlQ6bO1xpCTX2J1P9dPWLwlRkAeFiYzvnIw7z7nAbj7P+V5vKUOgS8OIjOAL
22UuDMssDjOhgB88iT5zuvPOR1e8F+YsMO9CeRAMbPGfk9D6YmadNbyqfX+t6fWKxSeUBGpJuIrI
eh9dmllbTGBiN2vLv+wMJjI4dSqzxdFMB6Haq5SRzNfx88Epf+O0pNbW4/DGXBP7o4GnV+u1TWQy
/7fvin1sK5V7SUPFd1K02DZ5QxexSxnClKrax5aeFpjn5vWO0a3Sh1e60V/6h4r7derFuDsVdhgf
TMPfzE/m2IDpN+D9u6Jzzw/YUTj0aj1JbkhoWNqnXNwnz2KFsogK2uoS+vTIXSAg0Hg/ecoU2sux
91T29bP5wG6hHGztR7SLurEgoPF+wG8I1HBPv6PhI+M+KrOxjYMWo5w4H/+aoyrFLWBT+DfxTK+K
laYATAdsGzY9Jgli0B/wV1xJvmnba6zPZtS+ROy7Z2pFE9KxZPPJvBoxmv759vM//IUtewRtZcPA
objxgqSBLWHnMBCkyumXLApsKwp1aGOB/c51CqupaqYoIQ0gzI7A/EwV5VQQXbk83Z7WigOZCQN+
ZFsvk20AvCTPp2d8aoEOCaAN39x1H5HbBMZnna9LqytCIeYS/doWd9EvEj7XyHS7imBRo4ZfOpa3
ODUJnRhotmGor7WZlFEgGq1gcPp103xm/K7IljHiD0CuaNoQy1Tm8+QXLhf4m1CnQc/eepA52yqa
vkhwAIoMCMgXU3KCZl37ArZ06gjg8kFNBX6cS+DxVK7mvkJL1vwZwn63HS5QJS/HIk+Co2A0zWbH
YWzTxZf2x7mHYRe5eVurCVH58S8QMzOkXjkkTVJ5eGnc06DPk6KrCV6h3Rvewsfo+5r5eDCaKUqJ
QqCFBX7Wo6KQJEG6TihWoxtaZcp3K4vrSdr1SG0uLXH544wRtOZFKVOs9tBmS0+w6/ZNTtLracOJ
nEWKP0E1cNzJXwmV5jI1xg0JmPoxxbXxa3mNBBMzVm4j7dKUTTzL6TBb6Z9PLtw3jyRaObBHuKUY
eq5FHSls9kbiFj7YGgUvXL81c2+O1FZqtMPFUs/tZWDVlkmDDn3dbfDfYDx+ngpPWs/CgAdeRNJi
ulNQL1V1Cee+G95FnGlPTdPtl25crNcfNp5vROHulKDRNh2Zncb6qtr8Ci9HLuSDmmzwyw3cLrA+
rjJ4gnS0Q4ypGGJU9kYbyCK6zYf0b8N50CAVWv/tvYkempaJ1X1d4Qj0SuvepBgKfVU31VLxEMft
b5Dwym4lgYR4rpDt4LMAwYafk2556AT8O75qlNroF7NLymdcJ+p7+zrIdwrVx1FMNXNTQ1mFNPvq
4LvZCPTtc1PI7dY5dCUTD7AQx1fUz5SfiQQzqDIS+887FxEGXrxv/tTxNyp+m41sNW3S5fj/AVgo
aow/Ymf0geejvl1vUaylZn6+dV1Jc73trBqJK0kHWQhJ255kOcpljHFvZYd5WZbdNVQ+nED+R+NE
CdF/lAk9VIgYPrqTcUAi32iaRb7tj/rTMXPbKZCJFjdBvWinHuCBZkgqtxPVCwrETX/sckTRtXUD
9SaFAIUsJraXuIeN0Do+avop55DiX0DcERcQGvmRlDedKEeTLAghgXwmBf8Dpas8rmfJEDM3Wqvd
HlMeORNGVeFMhnC3oqf1KEC5sNCuf5WvKbMwQ8kaiyIoKavSuqqnZlPycvKk5CPjIuu14NKxeuOc
PMWuzVdiz4G4u/xx4f++FzuAb+iBcNMzo0C6Xl/UsalrSJpFQIANMHe5zzwEvIoci1NdC7IaBK4F
Y/eLye0xevkoR4K6khw/iGxNoTuopCmltZtNvSbn4cwPjzK1QcqMszxR9okWPPRs08FVhqJi451H
Kg+/tJdnsvx0/9CcnF8Z2WoQVz+INffFqRzNwh8K4Ykhex/+JKTXsbNtdpqNJ4/X4OBI+13U6KN4
PgeeZDfNiYedfHcE0WUkQzImKyPvyAB3Yt1OXPkFtwjxUzmYYyXz9Mxh1Mhi1pV0fs3M7vgV/SDQ
P5oMughVURwmfQN75f5cvQY0b/Z+kt9GsmJCe/m1wlF5BcolfYLkILlSkp6AbpGZhKb2RR9ttSTH
Vj+MybMpinPkH8IKZndVWcPPVkvLxhyQ18wMDy/BwTM/Klf/xKTJQ2sMqEq2aclso7UBnymRhjQp
L1sqnOH6JL9hKrJXG186IAy2xOaJDwhNrpRPWJtmldNV1u9D3hCITsKeZ2eAkEU0R94PCjvpUsQW
MA0LIx/ZXvlmphQ5dDovyJzAtyTYixxvECwQuyKnMk8cStprGhVQhWCOjC4OmBe+R/iDCqRm6Loq
RpjtJHz48aFBHHWWiFw+PhYKVFLXJ4QnxolRLKK3IQP5E28iCSMaXXzuz6Jc9PWf6QfxlALq71pn
nBT2ZSHpOzIPbwFkHNfON3KLgaDDcvmYjTGJh0m6N7Cj9RUWw7wPLMdVIqvsWLcH9TRvHk2HAiC9
3HCwDi+5g93PU4F6KXYKKfIOYysxWtpNDSvZVt+L5+3rIqdS0zBqexNQN94t2yu0Wsx0XaRMnB/Q
Zb0WTLUJEiBW5X8+0EzFaPIUWTNOvj2dQLSFzTGZPoFc+TtQ5XZbXOD9Qh0Peh7nRH+O4ZW7okmY
MjVvy2PACHBEpvYMozZzvYQto6Mgpkmswy7uW3znRJqoCSwMhaJA1faA2dG46SLVTN1qGAND+Kac
xHRbiNr2TbOdlI+uxRVkzSJjpNmEzzQrZHyAfaqS5QoxtukzwdrFo4m6obe+FgAX2VdtcxH7T619
06LPV/vyzZ0HwKvZvWXhhlbD7T+ECk305uL46hr2ffcRmYbWzciLytzl8CpeqVYr1oJjv25ytOZU
qYN9aIcwSZ+wFT4+AOK+n50fefo9Ko+FJWiyYEh87evE/yX5RzbYTTOys5ZVUobqwNMh8IkS3dQT
dMChzhKIi83/fkvY1V6cqt56qIUiR/aasY/gIhaDIAGQdb1amNyHMvXj6Cb6l2VSL1TX0QgtFsDz
vo8jy1FhcZUDP6eM7c4f3NU7J3ukcB9iCSq33t1IUpZmQmmuEg+RqxaGQT3BE6uktel2LPkZUcAx
FzHcQz2kVR8D+iHkyY/jdtVzjF9UXyC1ZdRY4lEXiy3FcONA1PcT7afUTG7jEl5IFv4AQj7Ei/Zq
nIAIm3mWhm1kUfFaIntZpvqPEymtvmDNDOVz8kzBONaOdHkUiE7tCOi0DmucDdyjTXPhY+6JaNJa
ACLUOT+T41sWlYwP6LxChnI/jcZVVd2gGbUJOr3VYrx9KiNrQTl6QilMLbrpcGezxi60kGnbzSzS
jLh3auveK0are+C8XP80HOeciUHsFZoUWbDmyPsCSgiaZtqI+lo1ClIA4gRIesgCVCP02Bqeo1/Q
3seHPeWPCo2/FlFuB4ej/RAvX5ligwSGZkRESbv31Ik1Z04jN9RrCP/QxdxrBNmwmBvLYhxFzj7l
S7A3Rnc7tRoTaLyGaqY7FEjVYu+vpYGhfRU/qx4xe0EHG9BizSMB/Hn+BwO89jTrxic53mnE7ULt
z5/gbyN+VaRjKK5wnNnfZIn6jD6PGJMWrizgPYf9D25SDtwwDUpLvYf3IT7Sz+VMU/wCKkZ370u7
9V22MikphA7u28OvdGbtx4nOyQiePFYoiNZaesxuQ9FteQm7lQ89URbTCW5Yt5hhEFym4SpWPy+s
tcux5Lr4DPL6D5SeDu+TTH6AK6+3+2/g5L36fyaQj7dcatMcO2tOpTkTzSQeA2Nw4LAwk8jU5XhR
hMmWZjrcqittqEyHv4iGfgaQyoIHrxO/p16E2zMDlZPqKoLc+tccl+ghii6own2qGdhUMa860x0s
ar3DcbyD/1BCfbqckNF0Q9Se0W8CAJ3IENtxpdn/nuwjYbvmtWCP0zUbFoMALFjeQ38L00RdlGZ5
Vjm13H4ADoG9506KOeVL8zN8OOZiFKHK+Y3x+NESETZtrL9jfnrpoQjfH9E4sF6kCB9loYbmsdhO
J88GuvFyTEK+wxuSeSqg9OLSeTuDUW0zy6geT+Yg4249M6QUaP6zW6ycqaoBFcbsLjRPWVnfh+7N
uLTW7oFSzIAR75TviwD4uBjHrvtTfi/ksIs0fkhtWDZGTvVAT209C3nVmN0BfisJYhHFQ+HDLlA9
PPi3iQPeg6m0sgmotqgwSgiwnqlUaSikxouJnqUtV62ci0Gx7HnuiwEXbby0hzvXT/pPPW0+b5r2
VwhJiF2JGyAYMpn7x/oWlMKEicmnS8wDP8fFHRRtHn76jKAL2xqpUV+Wb6wluIqpMyiWTUleFlZa
dkoI3Fguqj5L1dj8WBDc5DPhOZ8pehfMhoP6POgd1d9o1axP8fs+CX13pwwAlGtnWS0g7iwd3T3P
n9EjYRu3INAlMsW1paLgO/GzwicmP+u1VIc2chs4Ybf1zjllrnGCV1d1fIBLxwMmm+INwSp4A0NQ
DmdnM0kErqKXqvQIk1eLvdKfLprEXFOUzRf3ziWjCSic7XOe1VaRrP3mv8QPF43MlQTuMHlOgDR/
GaCElnvue0c1hUdBLXEaxN8NOo1FTtsSungkkWFW84nKAMj/XweEx7lAwblhZa5zpmvTLJ086YBw
Rer9QzOF4GJMOB6cbJN6oprHfwFAdpAIj9MriKL95jY/255nQkgMm03U1c6IVoCbyyQzItnbPvsm
VP5iBMLETKa6TbdX4mZT20Kkg5dDhkp1ujN3t826j50FX/2Wu8SxCIOfwCle10itD0/NEwGtd3fa
T7yW/rdFMwTvAkeACYhJvKZDilaaiLRe0kG+6wRX4wCS0QqFokc3oSt77W+Zcfyi077//igZ4MzQ
+dvEJLJOGCm2Ic6hjukgNuLqxYv6xkHmITWWNAXqQcUEiePFYuvL7epHG6X0utbM+UVkt/ivZjwS
b6A85D8a6uvR1/1txqq4UeSKIaAzKJ7jOrDiwgYeuiAvmF+C0//jREXjQCUf9zKxHyEcBOPMR0/L
I8ehc1dV+NOFaOb53m8Zfpnb1A3KUrNbombQCww7zmVft+2U858Kk/x9zXh+0A4g5woWYavm+HTS
MqmD1LvlZ60kLvLw02oKcD4M4IHsfFQWj5tlfIIrC3BZC0BtcWFkSIKZrl2YRm5+GmaSHnz/EJK0
UCdJzFrIdyLOGRYCrRHlfhicRWPzk//Syt4Z8li9BdAo6e6wOBr4EUK2Npwq5vj1tp+Mxt1Dyu60
XCkQjfPg2Y7f2MtQypJut40iW6Zf1Ic6jJm/Nb9iym6wuVOn86jCjnT+uhBAHEQ6A5UvDiQffzPL
mycCVphFAsRxfrd/8f/09JQmHafyhirIrdHjDiS1Ah8DwdpKqVP7a/7AqWWd4g1IBOejS7k/dPXp
XwVReUD1m8Va7WtTkFer0TZyeWgR5r6rK5lKLa8JVlcpI6IQgPY556/QPBTdbh7WKvlQPTr77d78
niLZEek5qD8SmCZsx/ZzASAyp+2l3efrtRJqiRr45y4i9hlhru0MIgaOA9dC5lKMDKWWLKhKj/QL
sHCiz8iu8wUyaHiagCe3YGmrWIAsPGtwT7FUuGkadDOf+BaZiZnRN+RQkk8XeoS+nyrTyQBjgDAb
APvvQo3vbZSjeBH9N2e0Vn0Ce4RUMH6jvE4jOYRLxDT7ka6w7dYXnUTjzIHikOylw7guq4uqDQUO
85YdtCCARIDRpFtJD6nEnUQG/Z1anGvcQPU+2foAHhXrGN+KfFe9OMpM5CPIm5RZqexC/8a/K23d
wckUHFjnFruV+0QspX2Z9dPjQS6KHwsfVXVGbCJTS6QpJ8met/s81TD4n59FnWISoUwzLGVZvSaD
gEvvcS4lxBfvBJw8+rVSMoq2vuIP7NRIws8HvDHR4syx/5X/1AU2cQQAKHBD8JniWUFSZK0/AnvP
1TE5ehTCOah2EF8KPDBAIccz60wx+ZApjP8s3VRFe3VOgSfXxmiTySC6sQg3kVFJGUAnL3o95LWH
s1CLyDXOVTF9jRBEV41jN/NlPuSUiuFBemRmHy2ZDH/CcdQfe4gwNUzepydI7i6oG8UYOkzwLUnr
jQ4HBG8oRP14HVk0OxW1h9dYH90mjGDk0MqW5TiJfBhNDg7rjFbJ5AvdPlQDJ4eGtSDPkpwuJNqg
iUXGO61Upxojxz4RHMVU2OTTaL137FZo5nTixk+b92MJ69cXBO9GS0+80AFa17bIrr8GKcBLLBT3
yFdktMTHcSbGKAFWfkE1ld1jj4Fl7BtIuZ0I0VXkoZlQn2yExStY8T0DxnPrUt/wuC+Cps71I1E6
ym/rnYboR2fwWB2FvQzsLIRXUl9/P3VW2R0qxJcDgdw/+sWP0BBoeaDPOLXZ2r5gt2ghUfipeymi
TW0Yx3n3iOV1F2i1Estw5txOMN7HtO8aXWiY/0h2iUSNn0OLXdOZPsKjjLcjYkZyTH739Xdj4GST
NNdQr350VbweyNL3fr9NaoLYto4zxFEwiiF5DOEW6zLNnRScRoP+/Sbi/no3179yZF30Sa+oOPs7
KtbT87Vf4dS9eM44Be5rVbkiC4NZTEg6hPiO7OUevJ0RJlbv1y5btJD9kLE+HE3MlnBBBiGC3Nvb
iI5/hdVrjNJDcs1q7/Km3dyb7UcfmWhuKTfG3patlygrIzB+gqm1pQYkPiGqHA7qJIiZaU/0igDx
LTRztla/vZIEuUX87PLkBUtSdOvUuqCf6O4m75PgVlHjxYYXCt1kyKf6s8qhcapD32qLT+kzrQWY
vL2nd+oZ+IYLyJvepH04a/N63XAJ6Mx2naC/nMOskCJT8VhwpmxzjfQ/0Ku1LCmUKrZiUfDoNpcs
sOa2d8h6WfxSpnfdxrJiydZ2IAb9mmFIfIpkwia8yvkW+gJFWhzN6LitT682VWRT0WxeKmRFv/uE
4k/l9oNECx1ETWF7/x0ctZa5gvoyq9y4GVepuy+HS9b1Z3YuzeWZcpMCGeKI3MuBJ5d3293Q4sl7
BQ/fHSadYanIE4sLnAhiB4Ixa6KjWOrRoqZbBzr6/nKJKNXd+zU4yOxg3Fl7IMKZjtd/KVGqZXHN
i5dDBhN9TSwQwyrXBRCQy0HuJj4MS/Ww36aKwfGf0sYq3ROe9X8Mn8YjMUACGBB/Xf50ftXyBogt
/p488CMtz5lz5zEIu8CzGAP5gSD4gTXxwm9i5joCjQwNnulyZxCvBc39R9MMe4OwO/W0qOgZ965u
35ZoRsCNqRdXoR82H/5MSDJMI79lyD8UZx4L8OkvvaOkFeMo0VE3swSCmPZ+e6vRh7fgKWIhkjUf
Og7+qCyG36t3p5NyXdMg8C0HWilRdHKaiu1fg+EGZ2krPI/S8CkFSkeCa5C7H8nNPg5xoLb1sTFu
DHnAi7ydOnnyktw9xGGB3FDQ8LUnQMrXLZN7Q3Va4uUh0sRgtAMFBAe+oK4zVR72QLm3ZyEj2iD5
yfEdodKpcdZC3a4Xn5nYKU0ITNPBIzngB5DRejvfvprTRZ4/fmMZloOFY+KPnSh1u+n6OF1jTfb3
nJXZOnD4fdFm0pdzIAWCwll6FiDzH6odMLCwLqxruhQujN5JVBP1aj7B98nRh8FJEvLwTx3I7m7y
a+k8DnFRx+/NY8K3EjSzCWtQaj9KOgdkFtdMk0m2nnNyEm6ClAu77w6dq1HBanrHROcWh6TQ1Urc
9q0A+p9TAWC64YASsS6n19h7COVLV6uxI3/38StHx/CygQpI+GtjEvc5knG5MJjKN8rxSTcCJWB9
lJ+H02XKflfhT8D1luEQuCl/gg4re9sfLzf9NIczDWQo16KSH3caegtiFDo89/eKZqCwYo2LRI4W
bp55tGUDn3Tczfhaok5SVjD+18kFxavcsRUsSa8BOKqZMbtHZh3dKiSnlxJuJLCbNFzVmcvEgNmt
xFW2rf8F9A6jpKawoPeMqoZJ1FvLdgOGX/hsXHqEktY/IbKU4RGEXEnhK2iRRJpyMCcL9EnFqCB2
ZX6bqXE0KQ93MDhQo/RxUCIY64ZLRkbppKwsPzQRDoCw0sDyVwNAtneU3hvaoZ5aDcJrL41zyga0
cikUYAxtcp9bo6RlrMHlcXTcy77KdWjdE5xa/aUBUKLZLbk6May3/5mMD0BvouTC0RrXM7Sr1Dmt
9o0xkhqWAwXHnMb7AnpnZIcK+vOtJxHoZXIHN79mXLKSMILMBaj2GEO4NoxaTO224D25/hZJoT3l
jGtCBoPH2b8ohQRUz1naabgZmp1WmC53vEdRjUQqAgjeNa+LlAIcW1s/oCiY9FldIDbJH4Dasvgp
L4KT/kGz8Q58sZ8eNrZrNwlZnPhlsQqh4t2n3tv62nqVVHtb35GxaZyvF5KD5P5qy2Z7Xsu+yErQ
ZBSMQ13dnZgF/ajpUyGXL0C1md4npXF+up8/iCz0daR51OXEPD/h4OQaMJ86fYnchQ/zAUDx+8B9
UCcP5FNazYOMnlONGy2jmWXp4EcOAusIVKBznQQboNFT87HjqXv1JRJSAhQKeTPz1Baf6whidMZg
lfGM1mJqdJy36o1YrYuDFdHsNNcJdal8MYO5DMBlwkA/e5fOS8hcCUXiZc9e89IRBMjnj49BsYkj
CAtNueAcYuyKEu4/ak/0GCEleckn1LQPJ5bDcVxprj0JzyPuTCJ1s7aNAFC/R88t+GLcA9352Lnm
oNKs566QnHG+zGmKifCO5j9uvoNkjMArsQY89ZomkLBNBZDbsEPusTSagcpzoLNvRJUmdA5UWeGL
6sSt1sONooXvv4dmqOMfp9edFE/ibRGpcpJp+Q+EgqDFUrI7/qSnq/X9UH+Xz80ck3fnmf0n0cGq
Rm7czX/X9sY4ZfhUxSabXA1jVL9AYnAXDkLJiNAiymNx6IF2aThXDwzp27kPP6L4WmW+YC5ZNUzk
oIkCSLUrgag8PU4DnmdJZpbOzOI0vb+g/IngR6wuWC3vTA+tqmAKS6EcL4hMWlA19l+qHKESlbvH
kfLj6OouRoB8K83vUMsUPKznO2LEGmMahv0sO1rG8wOM/zCcfmqP+R/jttcCKxxUHpABqDqTMqYw
krBquTlRvjGeZg7Z1J8cIdh9MfJ+pT6OZ5z0PPbDOh11AWN+mECCHq13w5SUlNpS5Z6ne6qfOy4I
Ce/yiBrhC+5aU03s2jSyyIe5N5rV+UMbcdRBxto9ox95KuIWthIvEXOe7R2O4jOn2iYHS1yznlcm
stIReqU+Iop06Kfh59/7sKXQ7VjpVRhUsd3kDpP7WXB3JAp8nU7t/CN7U/mXnGd49X5HEAJlbRmZ
JjiDiAQAtDF7Sy32W5ltrfjkPHVevSy9hjIFQ9mNFen0oEpgrEnlKrYWmTkXoRX1TzhkCRBOUnn6
UkPAxv/1e8Hh07vf3N2kDQVRtICLNaR4p4wneHxBetU5jRZ+y4U6+lTJSD87FhEodaYYvuqAU/ba
wn73TZVr2bcEordWQHlZJhKJWqyq1Fsf0H2tGf3h4s8A73FxQtH9Qxpuv2qpP1RGVK/JpHXTPkdg
4/z0OVUWYp3jWzkd3ftWPIq0JFO1Vrm4eoVTRqTRtF80axHfbb4o8G57TL/IjH5CrA5DBkigSMBB
w/XQ4ugbD5md48cm3ShUeIkheMuMXaZEGGTNcZCcJdxPSUd1T1Z4jARD+CnLiQeOnZ0y8JXddeF2
iDxRVnEgAo64GRMRUHwxq7bfa/Xb8yobPDZEisbHRRUgnShq47Od464H/4swXuqmV2ATEBmkD/pA
1VFEBIrgxAGkuAC02N8cBdQEMWFfqrpTCI2H3bttUhgb6wq2U/CDeJDsyeHcH7Px412XC3koTSvb
tSnrpFJysI/PyPXf5icIs1FTeOOTj2g6TjJqJLrgjL2ZSmKFFpGXWE71iwmr/EzS/9VIfWwusDge
jbdioImezKiXreDT52/MBRZvFyzAYj03Lj8q3hQDoBV6uRekxZSJK/T5+CR2gDFTzKICO5jEfgni
c/sCOHzRKQORjfMSyhBReCfnp9aAOI/LNpWtbCbLU16Ghk4c4Bvj5x4e7vHF1SKOKEJL8nlI0w5l
qnEneNzZQY2hXnWxWJDbZoffL+CK08f2v4AC7eu86aGz8EGGR84INhmPBY9oNcDx4qx35Ga+N7OX
GXob0ZGD00h4+uN87S/msApGdqPe8pqg3/PMgL1CpolVqR2RSCghsxhJOl2w59xh+PAPj+JlRAWt
a9eECuz1dnAgzxHOP7nS3sCRKpAhuqbriGZIYZJuqKSVHz7FKjDpdJ6yOTRsSI7b2eEyweeSWFkM
AtwCGvZESvfGv0nMfW/OAKRxH7LusEPBCEaP3V9nxwwmgNEr3LjmAp5N3NJjbe2LQEFUUTw3/N9P
r7oVg6L3CGW55yCUeJIojCeJtRveujOw/bubQ0pCs5+l2FMoYS/5px5NX6rLW5mfy+9Uy7u8yWyC
vxEKCaXYnTXny9D0G/pxVptswGnUZ/5Ly1pWNOozZvgJRr5kg68zjn0GM3IHbKoKzaBpQ7rN4DZU
PnWDJmadPRGZ0izKJBl4kF3Ha09WDCEHIeH19d+g8cpHpCTs0Vl3TKEO47/pbQavCqgDjkCYlhK3
zF0fcGdHzsEUd3SSsCrvDheA6q1Qwb4xp1NMHTU2MP6XILxAmu3yX5xdNcDqN8plQGyBjyT79gqT
ixXOilzAMi7bIkr2hLIKVE/1b/w/pPVYOySGu2yIocx0nDIHxK19B3sl9AXU6iaJ45iRGo1bf2/u
Fc88NEoB/EDcJu1cPR7cTAwerpOBewIIYQjMHz+oD/9zR53H4bGBc14X9Lyp3dsIwquT7h6gt6/l
eg7+8NOMgwCw/ztz54nK9mUZrhJLWYZUGQStIC56pNJu9b9mOSfnEBcybEvEuN5QgdptICmhNX8M
Ljvv1LRIZVVsDRYnwo1ZSlFgr9ACLbDY4JogmnpDCfa6Hhsw9K3ghyN18W+mUGVcd3OkxxQQ3p4c
oMmkPETVuTf1YiW6SCra1r6XvMDTY9EOcGmNS+ZPOlPZAD+1UNe/h7qVLGfiY6jC5xQtkaLByJmO
le5+1inI6r5YA8143Vfpa+14PHoaYdMEZrjcGHU+03Ria4085EAWjjeV43VNAT9wm1AhckIcUys6
XDlK25rJcIVsij1zAqV/KnMlvOGREjSz28+19nkZupzcJc8yDGPgj7174+mN+ji22k7ipWi6kSUJ
qAsRbHyoNUosfpFUEKD/UWEJg5cwGY7eL8PY7gI1p89Yggt96Gg2inojvqOSKh3Lf703ERgruYUp
/d9yuPnZF2cihLRoy9Dc0A2eCkMtMQuvAsJ/uQJqKaJbVxCsvkhoWhjkdtsdtSJTg8nAeNTkdLj6
wA0NcNorZAx0Alh9Obj1g784unDDQ92NYkC4CGCDLvuaZSpROONCcJGF1u0QOpMoJq59MREM6/Vf
3tpQPAxTR8mqYNPTa3Rsocw+EisOxjUfmSo4r24RLkHxhKAv4v0cXDJLsMf/J6bPEhy/t/HdxyPP
d5U1WIJrpmxTptOU+ldWPAVScYRtb/f+nvxgyCcf35ySTMQDpoz+0tpyFetcZl3l+BnLp5eL0QX1
Gux5oDUuKmxXVQxEHDxbgpICp7C1grNHL0cX3iHbDpyObHFOzry4bW9DjvowUZt7ukAyoD/37vK2
frlWr0FXSc9uUR4JelkzVrB76cFDiq1eb2zocqsl/gZu/ilV0RGoUZ0qEnfLtSF4MRLb6XvsK355
RtRcsH1rPnqQ/Ynas9txIA9c03RBO5Iht5XKAcoApwi1gRi9kLMe5XoIUYRtnaEs+tkAH02Zx56l
rkSjJnLvxTXa3qy+wsgtX2+3yKEWB7nD8tHNoyW9u/EGH28mJOhv4xsXUdcJmo50HaexjdjeaQ5f
KNoKGXw9XrEyLsys7lIs3iUGXtj57MfJoBdoVXx2Ajm5WOP1Q9lgg6I38YrqwzVwygPfVlnA4TyL
BZAKWrlKOjcbSffW0dJyspAAhoUhNw/20Y85yY4wqn8AurWQLCdMug54x2kA+nle6hZC8KTJEVw3
x8BiY6UsHVeMDR4/eJvNzvbt2UHLTwqiROTy7Y9KcB3Sl9TcaVJ54VpVCm4xP3nk1gwV0WAyiF5m
sfhDrMGitZrXeSBMxyzQDBpK4HzpD6erR7RLuSViVJW/EovQ04rOWe5759k5m+7CR8Pe8v6WS01a
eZZsApANKprTx3NFCt2fe86PjldajGdTTvsKgvcwjEH6/0RQ22IsdBjrdryIRXvyAqsMbhM93zBb
/TI9tYsP3mJW7HtgWySqryAXc+oW1rQXq/DuZNeD83/U6AaAr9285Njdjas4N9XDvN6qfpatSxgW
LC8sSSAcXo3Wwrglpq7gLyD1DeK8B5K8MZrdceYLHKjzH13VDZncN0XdSb4nTimsG9sg5PrhmtcG
OGWoLJAnj3D0jIvEVD+V1TzzJo5+YPgPb547liJxdmvVazwqSrrQ+urRRcnXPcNigJM55xOGUxjT
jWxXc+PDlAoxv0QAIEruVQMRnnal1vSnd+PE/C3OFZrDxt05cxLfaCOuvrZleuMyNbDruNkx2kQV
MtR9of45s2MbEDIvisN0sAfTEoK5casCeuyeCUU6D53x+wBYeyqSGY2VbtK+BVwTe58xisWomIO2
ob8nzOUskfkQfdyHz72BGy6B1J6e6nGFMLXVyfUNLVahLw3tfTdwrhLPuZqmQeJdFNoKjeovc5je
CyhfnXqg+01o0aLgZdHweeGv5K2F4CJLyQ2SpC009S5cTIySDfj3qMOFLQ6rVZeVxQa4IrcluY63
YXqlYVanJ87ofeGPBwyE1NnWThWwCj2WnN4K0taRT7MycmvxEbefrKkmOwbynP3EDu880TO09hyl
AU38al42r0AwtDt8A8ccbjzddRcMV0irQw2iRkdXf/yTMeFx6qDlW3ujvKJO4+Vy58Q44gPCQJib
NeaQ0zASmfPEJdHrJPfsxs65FCdfRyf4c9RpB7czgsFc5KJIbJE7U3h/8yfge6O04a+QleIWe2SU
yZfZX/tXuH0vPeDsDsTrHuzaa1y2kqqSp6zMIby0Y91uSJkdNt9j9IbR7qkq4knb1Qi1qtna0bVx
xzAUNytFxhgJkT2RE45msaUA2JtEfJ0rT/6Les9EC2tSykNX6qg5RgoEL06jtSHy8Pqp3o1x2Awn
oJ5OIsF3IhmkAp06wlF8sakxdCN08Vmf4K3EgEG6zhS3MuXyCYAnpLjaJaiuQhKB2edLRerkmXiD
TO67Ut7S0p+qASjpStNQrMveumA0ndBiIfhm5g+H0JUGTslUP8T3l1UQsYXWbZAomJKh1tYvjpv5
BkTU/g87ZfzbMlgWU7ydtWzS/DWf4unXbHXRYEn0f/wd0JxFO2apfBWHSsUODUiilqNdY599KsBF
nr5AqMyD5dWTh51mKUUfu11CgQe/111r5sY3qUDlUAK3AIrbal70201TZ9wgtjL2YPPZoQfU8JhE
9Gjsu7okPKEmLpX3s3XDRIEVN8n97kf8gtKk5won4OIcslXCau+kMZsJRZeE6/lQmQ5YNPiy6rkI
FvBclLzb91paT7Rx5vz2NynVYiIPc/XD+9SChXYsrNGKqtm6uGxNupASfhtPAivk6q+If6QGZ806
7+bNvR9CekpaJU55IuFT8ecXScouqC9WnpOipKsXEaXxtK9HCHvU3WsJ5Nj3q8REJxgojlY+dxHZ
/iL4Hy2jcsE0ff1gATXt6+TWn0ryR+J1t6DZ1S5albFr/D6VxA13UqmNjwSgn8fX8o6PKCnbsMRI
urP14cqc4IRCLK+YqeShyWI/YZXXloWGk94FFbu+ibr0Zhyn4aVyEn5qC3Db7Z9tmyTLvrrNxe9i
2WxAtBWyA2sWsU4ebvCJ0O5ZXkzUpK/iZvGpWNA28jexG6NYXwWgJO7QJHij+LiGXybFJhLuqp7v
6o8GkmlH2OYsL5rzMnSUa43+/CS7xCH/g1703wXtrKgVwBoLbYKK7fN4l0T+UcPbGEFNTfepWkPM
ceWtuDz0ZsHk6FxvYENJSBmJKOtgPCeV2i1TVkMHKKL4gpLgc/VQptd8tUKY0gwrok4G15Y8wj3N
erofxZ6bKj82srJIc3KNphvON39lUFR2bofE1EEdi+uDHaB3juDTkv6P3n8vbP0deOTF2MvpFJHq
Rk28PEH1nTeYneYPmd+MqsreqKQ1mNxFDRtQw948Q5MN8ZaXzoUAAneB71SJAFpKD86oBmoIRBV2
oUDEBAm12nCBvp96kg6+KpqgizUCeR3TZYFH4CQYr3P9ptezjW0jnz9UOhnd4IaprFWy1F5cJtYz
28/d0MmOoVeHxWwzq/5w0uhkTdUTcCtrDgMJThJo0IJcIxz5PKpZabrdixZAMl+JqTxkOKq5gAyy
cf39DgVwn5X2ymVuj2xuq3HnieotidsLwalnNl/WEU3EeRlXIBAl1b5lghLgGKko6Tpw5ZmPdT2o
j/0qPk392VvAf1VK4dmA001yfnTur8XcLsabwuLMcOX74VKAJdj7PEMbLRvY2vPcFqmhW+vXNiVu
aR+YYQuC7vtgGsIqSAqnrn6oSYTkRrsdcjVLNN2NT+jB17mn7vTdV8GGCXTR7x0PtrmSser9m5e2
d1LnohHcUdD5bTNMmkuCBLYBfzLrE/Jw2ZtmZPo1wFZdZcRhOit/bMK4uNdtjHGFiKxQs+fh3IHI
ruU1r4bAZ/P2yLhirOOk75ujTlOvQPSObmBKezIluDXci/JCVVqkJ03PoNahf5MRNwHQYrR6m8ou
AoiMsJjnAAYetmLuRwbXZ7qkdR3uHcgPQlXmWguHAhhto0yrvIet2H32nYG0osPm1r+pXfEJi7XI
PzgeAjk+RHXTbznt6TftcOfphQ0gWdqC5gsfd98lT0QOO3+SCHuOJF6TOEOvyhZBcZqh2wfkvlaZ
bIpri9Nd2gbNidG7yl8yOa8MAt+hY4FAlNHBG6/kUjZJ+BzgZz3AmTON1/L94Pvjj7NpbXNARKBP
8lNnEm/jIBcRESYKkknNS8CTStSyRd5FgRCtgy+1ZNVwb4zIZYRHA+g8wz9RMCev1IsxyEgWerJr
Pb/qtCGCSj/UGD7Raq3Rsl0f6hExRcsZqXbBQKQhQ0W6UZX/cyxocHrFXEOQRhe6OS33IMWvPetM
GxR59DtUwqnJDwNLd2/aVUgZ1gY3noVW9g30t5fJgjucfKjOeGxJ/oCimQ41ntSN27J/D0919d2i
SIaydOTsuKVOQFtAavt+nkBUxUiJcRQ7zrLq/TRWVMJ/9Xua4IC0YyI0R1r6/oa53uX5vWMzteXX
cPSq4da7YSfdjcksTdjqPg2lMsP2p73SXnwQ8Uz3Df1PQFchHgQJscukMkN6a0GIRVhE0tNvVVX3
3Od1pXWA0luHwrz9WEvi/Ubeb0kgkl93SdVIcSpFlNPHlDIp5FkukFav2F30qXSI/2oYcaSpqfd5
iiCmPOuB357qfaOVzHqoo2xT0lcATG4O29/0NskIQ/qZMlb9dI3/0eqNXAFnIeRg7Llf77TNRJ3u
2xmAqx08HkVOWVGRQzHzsQJ1Ca3fe7R8tFWaEKfdBhiw8srBtfCqcnKLeSzWbcu0AwIm4+6vvILA
8B4M7WcJzhZxJ+KKgJ88G71z8jNC+hsjckRnjgxgqOpa7WJcxgijZXZFhl0xYp1uchJH1w6hneUT
n1/yv+LUETE1iJEXebA+6hIcgluTfP4YTwtj4ZHGPoCVwgyJu+D5+pNAhgIRu/t9Ehh4zTQt9zCs
xS2+D1o92KthNruntOx4VsFW5OkEzTHBE/44yykJ4XvwsywaOJ+ZuchTT99UgeLpz9Mp7xKKoF1K
4zXhaYLM12EL7EKqoYYWictWzzJaZViF0H40vUru6PKqOMQp6afEAcQ+/WUdi2AChZ4ZbrFQEy+i
XWVmpbjutHhNPaTUYgcYurqh4ExUUwLkyTLiSkKtB2tXzjSmGGbnAd4twrylBQ0a/YY8OOBAv6ca
uCWRTJcX4CQqBjJ7XogAp1bjaCMQIPNhH/oAE1ihDNe0+3OD3TZ98q0Y/L/8kqBXO7HOoCOpP7lu
dR2swOUVHUnoXeRh+oFQFB3q2qEa2WThyglVWBhI754JePckaarMB7gOUSrjK49aLmsR0W9TzNmo
oKxfK6IH5764zT4MIE9AGLgpxKWgUqxOyW6GxyucYUwEBhD69jlVz64ioqSFLwzMRT+bW3XXNVUN
s2V6NFCRuNsnU9l93GkGrfIApczRatuNyqsnM7kOHlNqH496mUCn7DvCcsWq73iok/ghcgjoJML5
932Vm9wJ4NJiM1BDObGkrnqfBVdpM7TAq6bP4TU1NrWuNEpImYCrI3OlKdLQuUMuf4jK0QsoKt+G
1oggaqSJs51g80vX56RrhP6vfAjFEbeO6q3hDkIAlYND8jQ3w+OJEkEKwY8ucGvxgFOQRKLOLDDP
IWtV/xysqiOe27J2uYJhEZXyGHuWRzyA1AJpnu3DFtlFGLiKj2vZS1qBIcWLM8zhyywB2Bll3Z0f
xoCEK41P5JFm/EFjkMgQZCCgnWOEvnA7NwRoqENbdUt0yvSQbA/GIBsLZ9LbzIsqXGy/qxXhtxZ+
DNNj/Y0bmMtpWduqPkp461er1uABg6te+0B+N7A2Hk9sKsoD6czwPxk6U23IFCSR5W3A1kOhRv+m
Bi4FI/0/bTabXytaWPL9aKmnr4ar/iKC0adLmkRllRx/CXklptVWAiq40XbG9pib1Do5Noktf8b4
Hb+qknXR7nr2VTYj21ikNsSo/z93n4kr8FOz5UN6oUd23IbhKw2mXc92ZWH6d0X1zGJN6JiHLlJn
Yr1JEDGBiWh6CCFxPf5D88JRUReOeaG5pMoRXhQpp3jcutYZCczHGqbjgSWn96zn2TKuUuVPBGc7
DLqj70pFF9i65ku6aY9Q05vfX8SaFXVCV0mM51qzq6CXzCldhsKS5pks8uiuOUlFj3dHXbz57PlG
xbKh05+IqeJuOs9gAFedRUlxmuPKB1ZdMcFDQv1Oh5KRQk+Kygl6JMfFe/bG6Ar/1SuP5I3qZ6YH
IiMpMtGeHPL7GoPWmkkJLMKIDHyPmy+6KgXNRfOkKnk2tjg1QXEh8wWv83uNFlIOW5xgXMIjPbbS
S2AmR5s2sh1xbhKzfr2dSpsPUSqKdwxpd8/g8+uvaNmCL7ugON1BdgC8TGhDpF6c8cEufSO7nmgU
ny6nPfLFuVlDZGJJrWNjFd+WN5DLJnuA4rCCnoEz27BzkNA3M5Ir5TpSRe2P+Cz1iAjM4Ujt8b/i
8QBeF+79GAuxGrSwpDjpSbcU8Y/MfNgH8eephPGYxZgtFgj7iGoWAIjg+FXZoHIGyOxmMw4XTg62
qUv+vubumWzXeGyQwocOdIVfmwfUqEcJFTN1UIlMufxTxpDTesQZp+sCRK+OLePY+LJhNTODPHwQ
zs2WajWYWTXjGykyMzcIhWLjJL03vSoLnY7bzMU2R5h3R4dtYqqkOo4ysF/lz0Xz8InEwfhC1JbJ
lCKLjeGgkCfd6v5s2gdY6Ze9dX/nkUDm/P65uXadHb5xi2kgthmiqt8tqk7SaNDt9kIh1xglcFu4
EK0ekXq6FXNhP/0of7y5fj8CiYC/9Xtf8xoFTD/2cCRTLeCXHeCo77SAUpgOzBQxnZr1GnXP3q3V
ATm6YX4zMt5f0JKM5AMJamHcmsl8g9zecZ4dW+UxPlGjnK7rxqxEMbqcp6bVIEFisHuEBrOyYMXg
nSwYLCzUwW4OlogssNl9U3rYvucNuBSQoHGHcfo/GVEfr41oyQ2bgIKuZANslqy16bPM7bNlo3op
6OzufvAfInZi51QJNoN4Z9hyyFu70ZodebecctuRFwnQogbr3SuFOPXySMV5sCADMMZMlV3bA7Ny
492L225fiOk+iuQfyDOfo4++G9zrfflcXZ7QHkVBTooDcgO0hEcxTThsER0ONjnoIEEYH5svQPKe
ciWiecEBPvJ7O0v9JFNyhY3rulvNmfGoAprcqYGp08wHNvx/Jtw1dBDd+tuAeIwp2iaa2aKreSPF
2bY+va0CKKZXC1OJxWLuDSup/UBcMfCdJO8qzsXSd1KpCRu7WFBPRss80VrNbWxCpLrlq+Wt2xva
SYXqA5jAyUzrYc9ZnaR7dWRVouX/Lnj3YkNo7VXOo9P2ydGbjQWRKebnJ1rWZ9k4zInmeaIHt9ey
u8WBROXsx1aNJIgiSCPhR/ldZ8YVY8qCdQ0UcywWZmD3iC1lFDF+skhfUCoGYoKn79rVaynuEPrN
eOvVMVqH2enUKBqYYpHLw+u0PLiCQhFYWmli4Oxg0Tg/dasKZXvlhHXqnEfNKr+pRb0jPueVZlzh
WcS3OHHt39sqR4reJ0xoUfxFd4OEZVzakTS02gYB9d0y79IrsA/nw6kUas3syjVHs3HJeqxd9fyd
tAfqL3mmXdWLFG9HtJiK9BRwlnC0ZRZ22289Lq27OcVzxJGQ9lvphRr04WiIRbsqOnnt4OUgSgYI
7rCAZtuQuZSbNXAb+2nrtCb3TcCIIeGdaXQONhf/C2/XXUiWn3YNEVeQ9R55Hc63CHvDBVlDntjD
xhXzyh84W4FqNuQyNv+Oh2BmYqfYxmtRebekV36yKRyBh1dh/TvW7Dn9f7jrGbQKjtkyQVR4QmTY
XYByvPrZlCeZFOo/VRayRP4DvG1m3zXaQwexrfEyFkYBwyHxEeAu2al27Q11bWLJIS7vc3CSyhpe
exZpcgTfOivrHQjgUuyY46JCX16XtMxNejwBkmUiuLVN1UGl6J2WJp/tsiB7XLqfQ9eZxG8VDB0g
W2pa2URAXnooJalMcrWhq3wmD0ybP7Zon5tMX8ULBcvqQDj0pNxgvUjnD19K5B1nIBKT02Ubt3gY
TypN1Pm5HGKVkR2Mh92LpmxacAVU6vJFOLfLFZD/ZOONTjGmpANJy3r/PZv/k+gzh6NGp3mndY+L
db4PEHsVvSDngafB3NpacoDS26ABPiaSjBIJCfOn3jWSDnp9NGnZ8yVfBjGjfM4eDqGhT1UItHib
FWedPKPoviTYySwTBYLjr4PYR/WfyQ5w8fxowAU4RzoFzIYvQI5P4iUcbb7wQL/Iv7zrzGole1Hk
SW/xvuhmhj2/3GK9jQOAUnZ2lPGo55lTKkCd3/OGgzrdtTBMetmNe5R4tWYFmIra8XtZajk9MkFj
x85QGpH+Csi6GZ0RRJPErl12E9pdyzbxx2ajt/jPH+2KAbV8CylUhAAPLPlEVMTn0tucv3bvDUDC
sRSp+197+j/N9ivuIOrveEtJQS7BQCHLjw9WVaISZbUTrY3eQDFv7Ms9WAGGFUvktQTPl/gVBXv+
+BBHNp1/2e8CXkjkCjIqXvw0UztdTKnHfzSrCwkBfYclGWTua13NuMLMSoIb/ty/SbLHMPIREkja
nP05q8XyOiufW5deGPl56UakgFbrxqBQ011LnUOdEZmJOPp8LsMvcIUYhvnwsn05Tr6gh0g70bmO
iWvJCDCZ+iQHp85zhaQVl3QW+4TNjrNGGMhzNO/lL60eakO7Pl0z+aHxaMt54g0un4V6bqA6ykFp
tkhTddH/sqZVfN1IeAY/5naNpgbM9Fb2+CfWl77ZrdayDt8zY++ZHdofD9R577LJooX7gL1T+iIg
Qm1iho+HbHYV37yDigzhWrsH2nJQUz190gnNkfRQCBKL9jb1ewUYkInqAdIOwzIp3+9EPq+a1eTt
msEc803xikldSVSHuL0nCkTYDWVn5/zrhvQ4wR7L7bqN9xH5SbMgKEibFr1AFt+dpUMB1QlyltdC
3BtfL6nI4CdAjkUS5CJWer6z+SyODSiDfOStN+loJOmlKia8nR6uHGixUoPX1XT2XiyGxsxkz/J2
lhpb2FMmiFqZRBfW99huVxhJR627fsXIUljudL3jmRvjy57DSkGeFdgoW39qOjCjA3u9LLfipwET
mhNHKijyXBk2M2O24d80d7zP/lSNzXdZgtTIewCwBWVYl1iAFT4Jl1Ij7xVsZ9+Fz0kCqkkMV+8v
eA1U4B6bujXely3vgu/SFqi/YDiyY2snCDb0mZ2x8W6TT0E5og581aArb7HWvh0d2QWInHGqOxZ2
ryB0/HxnH6LHcn7M4cyoAS0WfflT7UU+OmV22xCogS6qXpuf4Emw63lDTGBx4bo39yf0CHBwqDo1
IuqlQ30ERCzV6TfXspp4GxpXraX9BksjxGnC0Fs560cR/k+zGrA/dhodvnHoQ2Pv0keNXbPm4dpW
4chZXCYTb5RKYxyWxca/Qk4E5jap8zXrlC/FNMaRZjhZgMsZdg0foB0KBufA4p6ZkQ0a8sTtPh91
rXyy1KFuFm2hODK4kUhJkBruoHWwOAwuFpGwIkMpFocxYl5aP0vyij/gX/2z8SCY8MsDFhDAKvOW
o+ICt2O5ogsf+9lfYgsVlUa41aGDZvLjUxILTW9Abxg+OucoiuRIGrP8aEV6oPipnrAyxEQF1kvy
XAHOal9BgVJvAMBZUcJzQt6qVwC379V1wg6l+BtlpzeU0N1pUbwJe43t8dLxZwAdq1ffDuy5zxA+
RoKSf4PkFF2WQB35L6f7fmMeimDPHfryDHXrL9w94jv6ZtzyTbo2YoDPboOpd80lfH9SkZw+hju9
+Gw6qAb1Wkke3f9EmB4NGEtQBRjhbh816xXLhZ7ThGh8wloA73wKPHOrAaRRcv2/msxSOKucLzOL
L7Hg3y+lcuzSpGFpNehnwx/H7ICt1RCCXmd/W7pNCtOw4/7/WSAMsWZQLrbVfMoKKJwx3V3cGKhU
QRFkaIEZQio6qY3eL/sqhms6zZnsj4LZaNeP3whbTbW0TGS1I0NyYcBxpS4ATWA/Fw16jay28Z0A
xp21OEzvRS8hsg0rLrLXBi7Au5jXkyw7pBuPiIRdaosEF8of0tHk0CNaYRwZhmtNPcK8COPHs6v6
2Sz7epVhgjLBUz9+YCY77cEgVtpGrU+OYNnZfxmVqJae3r7+hwLJSo4vzehysaZAuGvoeUTtY1Pc
kNAgLQZLSE0b4v5shORg9Gh5SyxuvVaWmBya0ooW4xDlx2ugX3aIhPEoXtU9Bdu/X1HpBQkaeNjy
vq6E5w0H/3JsdcTC7mFkN30L3iwMvxsaMxePvKF8qa3fV2SCK5JkfrRyYXJ9o5DHArGR0W5VIXjd
z7GG1DZgjeRn3ALTmm+muH9eBGAujuZR9Y5IuBhifIiEgte7HCRS+qFvb3pN2a9LCcCpk/XYBeEU
NAl8mXyASwRbg7mXGfiayKtXcRshMQ/nl5hXDRaeBQvatdJ71PXByflGemBCChLUEW1VxJW2uEE6
SofRmwHcinhryCJx0HRU//qg66CtimRrI+uGKuI2M34/xl7pZ9JSbr8OlXi1cPtFS8RrNnE4b6en
dwmU7hEpG7hoLAAHxXcS8QeNaTfE9Ee7HjLpSkZtNW7Daq9RYiI9dk9f3LchEfMiVieEZQFB2UO9
/tcvojJhIdBO7WPZM/SqdprhU/XtACcMxA1h5S9844otXNXiPPG+UtWu6TzqQOXpdMfu3JsF62pM
5AdA2WdjssWPvS+RQlEPfCaeR/vf+arddgYLM/Shr2eucsMrDModHuz1BjpRVJrMNu23jo25zWX1
ary/XmLmrqGQpCRwAV0QnEU9rDR9bCuSSLIKkEkmEl2sWBOyjoD4IGbUNFC0YRCkydaH05bDSNkX
Q0C13u5PqxcLk1QapKM70hUANoAgA5vzB5U6ZIk1O4qVeBCrbHp82ciDeR3uyFtarD8KOQnd41kR
hdWIVj3t1D8m9k1xHFvMJaXs3QpslgGl+UO/0MqKNeS9IEV3/2zgGsvfkh6tLD6GW5qzANf/kew7
J76ns/TadDD6O2VDR/6QMfT/xsF/uIGQwJ3BadKfnLT2bHfGYRaLPug724LZHl8AsIMovGT9brOv
WMqFq9SO/EUCJHGGJFaK6qavQQ4/Cz0pvQM3IfxW+Q6kG1EJ/WIaEUA1YZPhJssDzSLcqLqU/tbw
LLhYbOarm41gX5h1FU+8wtyBSCTacnI4+Ag4QcRWcjMar+Lh+g7/RvTEd8jNyxl68dTFfLa1k2Tj
eoNyqRQH7+IfvXZYUi0m5TJXZO4vCEOA/ctevglc6M23XhP2zVt/ugrMIQrZSdKtPka3MbqTZyka
OuxOo09CHsfC2WOr5/0N/4aJxRS+mz3g2v5r9oXvzZKbZgz0/OF11D4SxfAsymDbqLxcmL1UlR3+
NsHMHrgedNXdG1JRV2Y4ov3HhCzjep8lWTByUKuMGLJvqsErfVtRYL606prh3Zn2UxWUUEu0OQi1
aiQ04V4M5g/KDtKAup9rRpu6PQGz/KLM0eXdcpt1DsLkMm3shIXN/17nU1GOF7F2qEzDJenID9xE
FHh/uwbZVj/dpD7thiWKMQdyn0P6Tjw7Vz1VSavEuZszDLuNOlQ6TQ1xfZu0KS2aYBWtBJBx2s0/
tvVklsmfFrBS6fMSlHMP9TDhsgZIigLODpRVJD398XeePkpwP9jBKmrEnTebmRRJ2BNfRQtWGA1D
wzLPfoobgKiMBwnGPgYkNQEeBUtO4b/M9lgV0n2dRV8BqaAVz4taEmcOk7kJkrGNew8LRQw4fBXp
P+elFYereUBqCG+npMCyZQWiBvf3hUCY4a6btJkUbBV5FhulFKYuaT7T54MaiZCIu+k30uwM1HrK
8d0jSV63BZj007tNWG3eA7hMSVHoOq9qdCSPpajX/Y+eIgUoCGKdrN898Vi6AAAaKFOJTX4fbL5A
oI3eq7PIcyRK/DwTBsclLTgn9/cL1taOznBboKgccm3YuVsaEFYcKIagZHtUu2OCxoM2KbbBpXIY
UI+97mE+QP9rKxOUUtDkEzc0n3Wyup3qPA1sZg7v4zLWZlC7CO0U8D8tCmkrh0q/C0E9K2LO5+p7
hauY3qFF0P3Q5rKiHxmGSQubPNwcbN8Yl+ao8depHSO2ISEHCucEbJk5L7JxoGel1L+XGdQoPYfP
0FSR3ih0TmGdf16GZjYSfIfZC7LR51iMLTaPaiWwFtqMFJQqmbFTqK0U7sxZ+6HPl5znZGcc2pSO
xZV6r9SrYkcS7zHa8O7P2AU2m75luFfjwzn+zXmpsNjnCFnGt6jcXtc8aCzog6yT+UMbFC/tfYu7
exvXpgJL375/xYix9s4e+Jf1X+/Zrn3p+g/oAcHRDGkEcKdwpvjj7+AYRps31p44VXlakswGvcCR
dKAVH3JAbunundhySCXp7qrxQB7AT1CYklixhAqk+KBSN33yIczBpD32e5PMTX1CzFJV43lS4LEb
d9eJRYSVY7iWMMCqeyKGrgfNzoIaYzKNGNFpFWgN8z1Go6aWPw1h2Yc0QGohQCzE1nWOCnytAqVR
dTHgXgsZk4OBWfpJKy2aXjsuF4otsmQwEZU4zDs0zgCCk3/6KC7ihLQc/MDeTYVcuEl5ZCjZq26F
dJDVnvwRFEDpszP48a+k/nfwDJmnm+BuWqS5hZXVHK+sbakuxxPTN8CQKjEcTAQzzujbVjLeQJDQ
pfS1lLyB7spWinot3HKUpx1/cjPM2tIVPtvu48Nsb0KKHvTOOfbNLjlUWUSy9u8BEsNXvHyw1TuJ
MB9lRzk+neebb5Y2hwreF9Cj6+zEW6d6a1na9I75fhaljL97suYT0pQdamVHTQbs6ku8fGJ7p5mG
a3JDuDn4PTFvfl/1Dl/kAsSGlV4wUh8oIan4g9Nh9Xnxksae1ef0A3NieTEnglyE7Jrroa8iJl3I
gwa4DRCq72ObFnXxnKNt9uskCAnk/C+ZO1CbyaAVE2lF+zB6PfGqtghRRopDhqO42k96EJ7+J+jI
OnkyHHd+Uo+o/z40zHU1UdPRl4tk0rwnFd5PlgzBAtTAdX/t2BedyQSZ3tPVWIYFP/W9XXb9mV61
mwqFomNz6LHnjz7SzDSX70Yt9fHvi7S8TnFKCN39rj58G1m9yhvxCt+Ggo6BL+H30pwMabt2iVAI
LbV69K8dRH6xtABm1Lp/y5fH8n+hcNVfU28vgOghN8vhW0ZZ/vyN0m5cX7rpreNBmkING4+efTnA
uleyiAaClXJcLktiio6QZpaPw5nCC197gAulWEhr0iuuF+fBI1er4zBUvTNk+S0Bt9R3xhbotWR3
pfB1tkMwRny9WTyByEVRt3SypOrg0ZuBz5tzKHeMwkOnkOcMqtcDcn2swe4qLFzbV2juleye6M5G
UjOpaTkgjR6+kjt4dCCqyPm+GKqwB52xEbk7GGiWB1AVHnYRnwylPEtQx/3qi4ovDUj60vZ6uKfP
t4/pZjpOTD7yDswbIEP9PTsi2iV8h09mJxjX859B8ihExgmpFWhz31ip36bmU9czeFXiyqIo2i8k
eB2VdW7D6khxtZVXhcEfhi9exlFbhOavuyWU3JYkrRvVkjDc+RUJrhVbWcYwUEQCpOgshQBOx8WH
SWvFccZ1MDyfMykvwm1mgbGyO9Z8iPT6KFy55XmFoZsgpFhNqjhLkD90yEjYUqanb3luH7pK6ktO
c+gCmA2f8RNQe2nVFkRNwO6oK6gbOGXZYU10Jq9EbEVwlTZmqkQt6dKHO7JcTka+5K7jX5p7BaNZ
6g47pIDFQ1/hRGYxZj+WH9wDvHG4fzqWH5DD7f7Cml1iYFa53vKxa11YMUbmnFf6uMa+XGNMprc7
BUIZTwQQrvk4WeiFayxx386fM8Q/QT91NBLmq/liZA96gE29Uud19p8D9z3ivrGl9/uFopzLbv/b
KrEwfADLT9rFmRAZSPmJUJdSGtfwqTwaUQDxS9bpSpWKPdK7sYPyUSQnu49Dfmlf2Y8+aQBBno8o
vOEJBPd9BrJj/9AHMy+HJ8VtoAw3fJh0DE/v5ZNBFN5Oyyu5ssXBa/3tEbjjENQubNasOr3Qjjq1
wIFw/afcOOIGewOCI5XeKsvtT1dfynLHbR+8YqgajOInWea9DMdu7pGHNRYUPlDhAg+iLj5j0l+P
75hv1qMFyoavRryIQJvs+fjFvR0bu+/RkHFZqsfqMjzSV0pnqgoxfCnJWEzakdtHdBbFZc0o5QqO
lckHpgxHT3PnSyHlDfvz0gdVcIiWO26OhQU7HeYKmxxASQNbYCO0NqYpLKWRqOoLE12EgxxRx2D9
IlsL4ql4ABv7c3Yvf83JMG+TmIAp6+aTHoSauPTgkZGRtP21J6lWtlQ222JOK4TiKTpbnpwOUmhR
lQMzdJ0wbOYE8RMzm7+qpBSO3t7B6lqTs6KT+YWGU/Nhe8PBsiNkdVeL8NgGlfTB9QEjhoN+Um89
yglUZVnieT4ezmXPXrHHVIwiWx8wf9dEwoRmJkfu7ftJK5IX8tdci8gujZOgGDHxgp04yakURXJu
EBg+UWXhIL5MHRqjp/fsqIYZCNGdnyTpFgv0x5Y3kHunB+ffReMy5/CSP5TgReXOkkZFnJoJRVGv
894z6uhAAke9vh9aaiemTzohOGfrBvaKZg6ZTkcJT2QAm9ByDUq1wg9lBebpfq4TJrbC/4kXGOj8
LN7+v1nSwS7KGKbgnVAGgyYIYdqBH1vi9uyh+CoTt+lfeOF9Vuvi+19GwwauIWjVMzFIT+JtGzdy
2l04H/xPUqjdhh7s2Uysio2D6lWHphWWHea5bZaBlJ2O3UWW+5BNKiUjn5w4lSyIzmn/dBRSv3s6
ZOiZkA9J92VUwD3A365PYEDwOG7JT1ja+jlBVKYzYKTTifTg06QASgUKpakLeIl+kUO4e8axGbm4
wH+9A3OoIWRuW5RfxImraPKqv2gsEae4WwteXNQuYR01RPX0D+2v7gI/09+NIlkP3E05Y1bP5BJT
eiagHGn9eR64Fc4ZKQSxIBCJq2xc5iMy5BBZ/JrFsEBr67QTTvlhH0e6O9JCKW74Vk0buhBD4WQ+
KY/r8qbfrgo5u8PDitZiQcwtwtpnEGLiRn5h3CCC+e7QRcuFKnFLG6BvXxacfZVbITfFfz0enOVy
pgwPPHu8t3XzDQ3bsdSHyzdw6r+X7pYIfu3K8EOoJMbB+FVDUKSm3IdkL/XJsZtBg+ws0id9ptjY
1AoPT27X/2YGTiyhwCGCQGa7qANjbNhhVeMMchcF26ikSEc7lAqHsFb1ygFYMbJaRuL5bBFWYS2o
jw/cKVYhbiscbQbJDZr5uc9EchtSlJPHj4zXLnJaKo09YG1zI7i8/D9v4PPBQ44RhE8Qfg0x3hbx
V+SNoWrDve1uxPFf/lYLO0cZtIvcexbvmuzU0U67bvixzMQAYDHDp+qumd1698iU+AnyHU4BSiC9
Ijr285VgwrigwRNCCxRVhLdZ2hEr35cpp3EkYrW9fxVLsZgytFkvaXL9mXQFmwSULPeF1Jq8Sbid
XsH1KwD3zaKs3LQGyNnyy3XGfPvJr0qNyIqmEc8hfnv069vzccQCxaw6en8fo1sTeyqL0U0RiDs0
8VzpDcmN4mPoZ2UC7YsJzZ+EAAUT2B5Du8522YVg8vZaQSGg+ELhKseGwWiSopHA3Fs01yg17uX0
vLrx5RJofJr7Zz7QhNKJmzk84+T+b0UPyuz3TitFvN1hpk86qmv4L3J3fEvyL8/L/pcY8wonnGul
HB8hVSJbp0K99Nsmwxe/ss34zFDZQdaB5P1cFw6n+24g+AOtjDvJjv9HxHvk9yE6pQXZq/sOg0wS
dliCSOUe+AHHVAD4vLOMWo/5fxWIrMRKye8UB4ozntwZdf8yX4ApQ0a2TLBfIk1v1/uyOWpWOmFs
mD/4w79fDpjvGNgcMMhJarWHTz5TXJYRgUOpmWAqkoZXTHQsika27agi938w52iKqqe90S3kX2Kv
cGGkXb5nT8mjOb88ZvEglz/v8mFbLigKgKTiUzSTWL5Xk6BWfiPdzJGN9J5TQvP8GU0/7rWiCvGA
fx4TMY0sAa6iQm7JUsy2dk7HNi3O7qCStcM7eLpFrVjZPrxF/9fToK764DQRMFXt2zHIfZjExc1Y
TMGs66KQcM+3D7vSjvvAj+7aFYTw+T/e7tBYGe3M8gQECxijLja4mSoASPOBDIs6zkQGOj14T9Ye
G5pTluimhgqYXFw4xEkFIs0L8QTZ6IO72ZFsfFjhJhdt/RppJSpa4S8JPoaL0/bz4U5ugCptvcBN
/g/igwDDZ+DakGlaQbYxOlqY0MM5rYO+e55vpry90ixtWQjHGyrT4dVMC3Fnx1S8BOsXb7L4YRpT
bxaFj5420nXH9AOe+EZUhgZVwJGzH1wB8IGcwnmB6NPDfYA554dRBtp4ikJDsBsaCNJOl7kiUBc9
REbmCBCCr26iREfG5XyZoMxTxO81pPZpARP3bkB/I9eAvc/FW3lI1BAJUTDYONP5QSesjbzzkiXd
bTqkIxv/Q32X2xixy+w/6x64LdsWceztOCTTbD1BRdkHzxtqzaExdeUMuhiqWHjwrOlDJJhlgwwG
fW0SFAhAl9bIyje7/NW0IClWdrYwBTqG1h9raSKrPgyPV2bkXjALT8HLrwqWVB6Mj9co9jV9WpVP
i48JUFV/29yfCUdXIEgk1Q41a519zj8pN6t22UhcxevzHwYCnKWcljs+Qkrrq77Q5nU1KR6ZCr5c
zE7nym/LBAl15ZwQr8eETVLHrTVYAjpPvjq7QtaIGW8khdXk8y05wfWcVZ3w0G06T49eVdeEdnhC
WsnWt0yb921kleNZXoQMFP8TtjvnbVDMngkqR3gKaiyO5CNWCFR0pmuw3ZrOjz02yi+nnHlRKAi8
AtkJzy1dFb2v+I0VSJui7HQsXHzoA14QvZD8Z1kMzfj1plchikCTVePVi3XNfaLp21XXhZJSI7/E
WaNt30Hdl1yNLYmeqDOWZMJV/Io1o/atzmt4p8EWOruqZkTHMNtQGTZHhZPD0prYq2t047qQpXeq
/s8K69es9VA+0tXN2BraJ8A57hRkGQcVWnRGeTmc/L2o0PdECrdevLCpVm2/EammFGhQl9qJncs3
v4K5fL2IBhf+kNsdXXf3pHln+rSyrwC2CCLATM1LR0SZ54zX4QN8ySKUnhoVKH4VtM3r24aZwC4R
WFVifkmzABIMnKEB6bOlTq2QxO1oLYGWmRccLLVIMJUOva+AwEDn73MQDqxVbJL0YovGPDsQ/fTh
hRS74gWxY3RBWmaoYv6Aa3gZiU/bLBe6jZJFqrZhvm97Z7pdVnJwTDEGPVWpErc+tsrRBkM02uzR
OOJdeYPXrjWzMQMtwaHbORJUlsDynYlaIfBpmt3Tk1LoyQ3AfxwRLDPgRGFtYdROrStJZzXEx4wi
QYjDn7YVSh8p4VOPI7gl3Dbd2Y5zhrQ1bqyemIHcUu+un/XJ1qyz/NSOzWASYEcjhfCEdNa4Ue72
jtReizkuSYe5pT2Q0go9xpuWZF67oIawntypkM4u5oE3lbbebQL+EtnAv4tikpha3m1dWvhlzY+i
BOei5EaEaaoaogWGUJ7Aig+OWA3LcjXtsHMRT40+D/G5zEBd+cGTOBTxI0Bm4fa61EersXrs8yun
xJBfJSpUXQ/od1anYwoORX7Wm6vGqWsD5mHHgkhoiv6C7eTiSrBsXYDfjgrqcjdH2VlW8RjkeypC
6Je+gR5IwCNL6w23dKi7FfP7/HjFO6I5lgTfTzlkdNPm3223sNbW23H+gRGckcBeBCE0BSCKh8vT
nv83pkWMqapSc/8JVq963WGs3DWqr/tpkljXqG/s21PytIS8GOfmT3c0beEfK7grUVZl3T6WTo/W
pQGVddCbx0ldyYmoxpgbQlmR1R+/nJE1bmSQpEV3yEnzFH+Gw03QzCsFa0CjMd3ukmdWTrne+zuO
Pn/MkvEBfzbzhLQWa74pEJDgbUdGbaw7grzu88t2+/1LZYezpY283bbKEhB14hKnYtl1rOFVyPF4
r5fjxG68W4etEw0aKxA2cKPee/FOkFF6WvgS3tm6dWX526JUFPSmXVWS9lvjgYB9SufueaCnoIM7
mbUcOPiXDEoirezwI65NmnuUO3HtNEXxSWKQi603SiZr6CSJPYC+mZkR29FrogFYWqvgcqfGg/2x
SvTUVVFG9ffBWH5T+dQp2Cml6ArJB7nNJETwB0BVlB4Oj6TzygVHL/PCW5mO4g+hSrm62BBQl5TW
mgCr2KF3x4Yn46ToICh4VGR827K7fzSkLgnXgPCpleKPX4Bu4L0Yb4kpLRljhWHA5EkluSVR0Thc
/qhZfn4mWgpNKdt6dtITEOOAUzTR2JbGcyMHyGpZR1fwyT7JmElcFfOBlaHEgluxv1gdJTaNPdW8
rhBlbOd8xx0twRHU1MXdzKR5w71o0+XKi6TCsMz5K3gr1ZJx3zX+VbSnzsK/S99FSO9WrUriPBzB
P+4WMK8JN0z4M61vy/U48Kf3xYKA/7LxZG9gHqMgEmrVGzR4ENEOBiQgzTYkEoSvpmh7GC966Pj4
FT9Dvp86sV4D5GqrO0mceYhc0G4+lj/x1KiWw1q8SoGM2S88nz18AkywCuqLbLuVfXf9fT9+DmHD
xlxsemKdvO3IwSpiddn2CR3QdIgQK/WGn0IAXxw0qBHlPgsIU+LFMQITjrLmBDIIfCVF1xyYYqN3
PSZFw6zU8BmNBfvREnU/ApyKGMPk8MJCNg/Asf8YrH4Eg2NRCIPcBBPCh5lOmG/7CDM35eUFrnXP
Abt4tLK8PidXdbacsuvk52bCXtAhujb69FnzfjITzMP/i87HNLNqt80SIzCO+AIapr8qIENqaske
5iABXJdJ3l9pfSjT5wvqXU0gnDTSDhOB6VTSsq7/JyfZaGBkSsjVo058S4mCcFqLns1dLR8OJD7d
H/0hT8mBc50wBvwvuHR7LBF2AdFIEjO+6ADPmEVdIyTynXswk+E6LIKl4skh424TR+YUlZuHtlFl
ssZpbXNrq6KU5w4AnSZpjrBWo6qnjLLMn4bUevCMr93m5aOj0KDgL0V4a+lVomroO76eJWuIJTY+
pVNfhpMb8tZ63Ak5ogIX49i2NkMz0nugJAvOthR1lSMpg8qfhmyVnbAyzi5ltP2qcd/8bDpd6X90
2RpMtmT7xIwUc6FpnkT0BNd2Q+H8vYrAn+4SdJiAzntyjr5jYBZseKD4l9Osin9jfXxY+TZRZj8I
/FqvagW6Tx9yYgBmUExoX2AD5uvPsIW4UixD/mGjtU3CuhbGaMgBimnuniydBplLmDn9xS9+rvn4
b9ymUxjH+kJeMgKRH4YQ5n4QD6nZpr9uwhjOFqsc3P8Qel+D4WnlVCvS9gg85GHqnDBC/Wx8EMLa
deUMqTHObcy9gBnNb0NB4lmaZWqyOV1+bWNCm67q3KHdJaVUPGNFTVkR+ZXPAgnEyz2Ean439gks
XpoQH55J1TNNV+n6Wamnjkp2y/RRIsU9hdD4bDgUo4ZCjwnAi979sGbhyqK6KlP3k/tRWIp4ZqV9
I/dhzr9ocFo8znRq6dG9HxR54aUeh1Nx8b9U3jmqUlhaur6/PWrqEOsUxDZb/84w80pEkeSCnIhD
ILUKqn5A0cY9JmKNdLu1w/dir95sV7vchE9WhlO91NMQ/uthj3Byq5lxngzwBuNkfWDonSmk/ywI
RhMxjTHzslqLXPR9JTz4GUPtm2KxFHxM52JErJiILtc6aldBLBAKTqBMG7HmVbdMLq8RWRNWQ7/G
KIEr2VpWen8dfz72WW7l/OO3xjIuSdc0GWSUYwe+XO6NPluG6IwIWjTf7ecvV0fW3qsqxZiNdOUn
kY8mWw9s7XnN6XSMU/q+wQzufPGUAnRqWPGkZqddzH3D9XIMIn0YcJdU67lAEUxVsizHHsD/aO6S
bmAtRiwIniTr7gNIPfB3OxWgTkAsVas3K4jE6do5AMsGbYB9NVXawOLkWXWawN4XR2VYmH2Q0vBO
8xTlDDyauekS2UmW7xaCzSjouk0QDpT0u1iBlhkM5LYRwkjE250r4ZNnE6iExwBuo7o85uMhNy9y
D0nDo86c0d41XF2j8+EIPzfscIAKbuSkBm/4CNSffXoG8Ra1tFAffGBq62vEY9Y0gN2wQ1aq8OD3
E4U5adEsifUel1gVzPWJApQGGVuBqZ9SiRrmlC2oTeA/vqhOzaRzniNgUkVgIiLNv/qr/mCbtijI
gwT2a4oW1R5OjbF5uP3OokxlwlI+9NmhRP/y+kg9qkf7WGiDnjlaieckqWxrm8HmELJQHW76ecpo
ou6Me9H29nBz9hpTny2Dr4GaFveDJFMSmY2RlMkgnqso+lNojgy8siu4g7vBvdkU1QuMCfjB3Wvi
+MSIpGxUe1AibOoApXbT8h5Num0tnssCizwAmbMobp/DEka0zAq+TrbXZRXD9+KyHZ7gP4LL9Kzm
o8d8bDZeD025DBU5MP2/f4wbhck3wvKEpCxiv3dRK2c5u1s7MTUPEwuIV+oUxwdCFoioXxMEi30Q
66cHy1+LUcDJHC9Lt3LJQJroFdg6ItYbDeFIPWKxiPF8MW2ekRgOiXYSPHkqQqg8kPjv5sS0oU4A
tqLwN8kO7xnOYDebuHWJfvapviUUSJLB+IEujLPXR/NZriGY5/W4DOGRxIp7Rj95vQg+PktkfQ/E
DdWv5pYNQTfV86PC5IHjPyTBuoLdbjgmr91hYMdpD3kUd+GvwfCj+kQSrLbgtJ8wAuOZ66vB9SJA
/70YaBEl61L9MwRo1fyxvPS6t6y6LC+LC/M3l53WZRWL45gSUzKbk4pAv8o4REUsM3jYqh46Mkx5
EIUyvYBhc90xxdFQ3wGhRnFVDUOOI9qIyHQ1a3x8wowocYz5BhFTaNB9HIK+rEI/XdUftcMWY1ST
sZfRdf/bcNF/kSnCNmcF//eUDb74OaxMsqo1vugTSzriE8OMSNaZ7EgS1LBJYowxTM5PNJ4MX99H
jbe78gVBj/TYm7oKUYLKSseKirf11Z58UUXRlX8ChGac7lZ3qivCYhXNQpXCCNUgrVJN9AA0Dqae
BZRWfSkPzlG29ePYQjg7i9dKzTmzCh8uvx23CgONBikiTrLOOfqhZGBFLjAGnt0Cd4HKmEHXemZr
u5Yl1mAaHnD57bioIGB0LPhhyhwPa8tj09Z3bIUFB8TNOR1/RK4uWMG67YAPhac/rcc0+oYnGx+A
q31U/RpwDynAVmMYR0EzX/IY3divUclnUsXKViKyfkYlWPj61sLriS5Uu4XRcBi51w62mJA81dJR
UoO93WKUTzmKkuZo/8Q264c3GZAzJtnvl1m7i+SKZA8joH99hEx2OuMMj7gCheJGlQXHEXqmwaHl
y8gR+Zt7sYRtdw5PEcXgErfvcNXuuw5BPHrgLUbXQUFYyM14J2IP4DAazLn88eNV9FbjBHD0a0OE
lSTyKqFqAVDm+AAfWXGRy6bZik9ya9CYUmhuS3Wh1Me43DCIMXd9Bwgvgyvln4sR5RGp1erbRSZI
/YO56/2pnVGQOy3NgxbG46BYRAq21LB7L04Gpb52CIM8NuLFQeQrfz0v5iZUCzdUEAbk6jfjoXGq
LtB4QrYcopJPas9ry5ZCR+1ok2ya2wGAgSrGiLInx6oU39zPwHXMCMxU3cE5qGv37+fqtIPelJMf
y6MZVxWunBRQqYz56WQAmHEJkMb9X8rjkY7s1t2/YZ2l/xhRK4+Ndmhn4hJWwtDiJaPumS5NCUlv
wr8PnEP0wfiowpgQkzV340kBLZ2Qvn/9bDF4v4lf+rIftxJQtOCcxChY0/pNN+hiXfJEpxl9j31D
0ccdH3+Fjzo6oJI1jUhViydf6EZaBM0p3e8EaNpUKrdOJE00TCjVfj8mqBZtstq6BX9WzokN+ClS
uZ3dPm/S8y3JMzn30tyrgJtusPfN6oK355gTgdgRWKgulmcqRyx9KIdOdtC2/YkPDFQ6DrIHg9QS
8Z/EY02vD/h1E/OrHzwrj4ixIRaSofBdFqAbbgWkTkdj64Qh9EjoUm7Vn9Iqxw0R3fmu70P49KW6
S4t9KRAxH6dCuPl1/S8hnwKYPgvqnhaYSOtgBoHEUo4v/VIeDJMH2ynZTkQbdc62inYnGWDspbRz
i6bYy9FqjbPNXuQMJ2AVL/EQyRMWlLI8gRtPN82Qfg67/t4ikS1txEIhcnEUDikb16gxNyyz+ZmY
hSLIvj5GmZB1Aoy7DgWE8aCAE4wn5grI7Io6hqm4lpw6yCnDuEciMAAJibTY0CHifBrnPGsIOaay
Mgqx3gOiG937aQTiPun0dThbVCMeOjdExXGL0yvGoXzAyjVUGl+w6JN6jxbUjlrqIJaXU96Nf7Dw
JB47WZAHnjvbVRX7hJCcr3UZ78PStsU0a6iQ1gVIHcZRX8pyOVQC5w3trYeUXqa3rb+xsqNrBL2u
qgcbZD7/6GSilSATQu4xHFp3ClCIY9nGFnq//o8ZFt9wb4gWKg6LJ3DCyaHKHdYPbUE4On1EDcc4
U3+EDHAcSQmSCslN1SUhP0s7iU8I8NvNq22MItkAkWhyiyaeSa6TzjWRDi+wJERzpeeUt6TmSsuj
wqoTyIbdv/my0azk6fsY8t4L6SE/gP/PsgQVf60CX6XpzI53RMzoN5q5L+akVc86Khntuf7vEnwP
im+AMo5pgv2x/aibwcyIIx4MkI+BZRrJ2wFublU5R5Z5s3F3duPc94GCG2dhy21nk2EmFSJgRsnE
4+rNdxBPHJ/FFfLhMVDxLyML/4wvLt5rA7tD4aOf4p94c0Tmquu70S9onSkHlJeraFR7Rt/y58hc
TlUfVt8H8T7xtLwUir88A7kqRDVQnGH0SD0AcX3TfNsiywur2OgoLFFrpIOMZDynSL1Gq88vhCFV
93u3ZTug12v4+D6Cw9AgRVeiLj82nODRRlffLbJbvH1xc2ZxR8y5PXkcQpr5O71YbpR6JVXI3VF7
4O6VUPFskJoAPdDWu8aEmyP+JYpBLaVfklSbYs6O7fTDUO8qa5CU0OlGukgGAupQ86iYrcl9M2/w
n9qk8UpVNVRnTWfyZWFYMgSYqMbS/OL09n6aHg/yytSxg68xobHsZ++Ac4Wzsqw/e+HgHAiZHbdm
E1Vnu7w0jNsoaMJieiV3MTlw9patuXZ2QqNdH6dBvv6YqeLAjn9jcq3WXa3vMB18tGDFJueLq65M
8D9LNa+20v/zLcJp8Br8oSSX+ZvSqhPB9zNKqL6u2w+q/BoiJRrKznQV1B11YeJ9/bZfYj56cfW0
D0tdM+4N1IGA1teXZnij3f5wzH7n8xNCA2uL3dyZn+L0ZsPG8XuoTD054HEs59Yjj9ZPhmEBGP9y
rPz/zrrvNTqLgkHMxU2z1GuAWX/Lw7rBhZNvLTdZRf1NTNIL4Oo5oOvV0Q1W1koTDBllJ1ItRKEV
wki2GLETdW9ESxQsui16xpox6HTSvKtzBFLz8qUVaA6/ckH/sz1XPR4c6c/ShYI50GXd9E9X//vt
UHqkMKTulKLhVediyGF1f1tlhPdLAL594LTK19azXYLDQ0gb7DFTEKxuL30+vJC6CRcRB/+fDGSe
KpjSEL8slXCTVX65fkTSE9qs/TVmeEx4mE2OgZ6DFXlU5Z1nLFiyNSSK6zi+uBmsL/8L2dQZe/KU
6//4OWct7OMHitaPg/B4yX7OLSjHhO1WJAp16lqe7jd4ZK49jta0KcV9MqTi6JtgrOHKyiWk9SVQ
pN7X8vTTtltFbauM3ckbj0fCMyQBiJapceRIX+zDY+lLy51lcge5zmALGaRu6L8/zs3nIPKJ0MAh
S17IfaD1ySAubvkbkYYIUVJJwgSenqpyB9/oOPfSP5oh88KYfz4iE4a5tYf0WG/5/TV9de2Qg1Lu
ZkoT4fupQq4SD1m5rVe4gnx6szHgNkH5yN0w7ip9TCeQgUCe/PiuC8KIvIkKAkt1ggRZNNZcp15G
o8MUSudj6bkgbDhDckeyV4b+SpU03OydLIP7E8yTzJ/Q3dJIodIskmJn7QQUNR/C03s6iSpOpHrP
XbLXznq1/CyPfsRx+iHtKlrTq3CmB5cZOdyYK/oYXzCxegJlYTrK8wuET9fDJ2R9IgOHBLhJ0Ptq
04hZiZdaurCvS/Q03YHjyWPxr5HgG2HyzXM3RPWm/kTFJ+drP/GBHz/dCLQO0RndKMrrmxS4TfSJ
LqTaHBKaGL/8ppxlzoh2ows9RCwcHrGA3XSP/RYpYB4pE9qH/Ae0EKuG7qCsPdTSmeHBKNT6M7dE
lqSQdPi9vYhpE+FPHyCzG7l5AlHWQqbSrBGj7u0CuzgUYtkHA3OujxoQE8wzvtlaML4Mn2dwKAxS
KYUWl3ziWAKSaCN9eGbqI4GUDeTE/eUbUYZFMdWaL8mR8dmaZr2jCz6Rdw25QY96Mpfs+H8dsqkb
w9zNQbdlLlrm/uVBKzxF6ynX7Tbhzd7krbL94mzeokBllUTqsREw0fW4s+PhBbkRYizrAUDkQBI1
xxxpAS2g2F7ZrINZ8JL06I+XM/aBeEtjMtgxTM5mEErsTVfv1ODNBbvX6tSLkhx770GMAug0F485
BamQrlFMIwla1c1w1cyIYmxxkJa3Vk9+g19/IBbIL2gZGiIJTvSwOy0s60yNjF7TKoURuwofrcjS
X3IRWIGFEvvi261t2QzhciYkpaE25+5V7MXT32f3JcpAUfdJepaeZllMu89eRSuM1Eu12W3FKqTX
iH2mjpxiZ7bc11c+7BLkSqk3k3y1Jh1ZsS44ZJuLKAxh/Dxnbbo9V+9/OagVYE5aYsC7dugqvDIL
N7argt26c8pgHmrptIgfJVsWx+r9BWIoC+yYwr/e9rLAMsSybtLRccMtBPq3sIV9p/6CY8LILo1z
xWltsZiID4rGid1bz5f/k+vpYsrNmDfEgfUmearNVinjGjC7Onvjgns+RViXKybeh/jBnguB23sr
03N8jaTXT2aT3i2RPBNc8MfCjzbqm4BV0EZpGbfGkhmCxEnCzQagm5/Dncbvz4L4Gdux3OIkpjrw
dxjVPUd0E3C5U098Ml6t/FyL5vOGW2Ktb/M+R8oMGRflEw0kHllvdw7kvFO7J4eLz/P1dfZTXWnb
25ixjcMedD4vpEzVGB7XIZaYmg5NIeN9vsIpR+2L1vsAVBrxBDolD7UFRN8feQwXLUYiIkt3MQst
RW6X08YX9172ST8VGRDTZmwiXfR4y3FjktVeV6xaVdpY4KqN2wyuxjii1KD0wwJaLwgMrau0/5XW
r3HYFxF1boe/O1TlswJwGQHeCZyyJSVffYDS8oYgZRtcxy6REwy7ipdBKOYGYogIG7tJQkNpypG6
j/W/qWcyFIIeYM8QnYqij35LsT0Xprtvj4PQ4rNRYlky6nDz6fHnZw/MFrcSczgjeEUDg5LaId3p
tYUXlwZFDjATXnrQngSTReu0KUteqZTGAAkSISeZz5xmYkdsWx+MbnvXzcaq0N5vr/xp+5dTLIqt
B/qx6HKrQvdCTZc/eMsn5A083OoENCZWtdrUBSJK+n+ve11g+W1Y57/gNZL1kQfluexryRb1FUqt
6X/s83zjiudP5Y7a52Sy/UoY353i3KtrX/Fiv4bex8Ml0j0LsYdi5WSr5wJwdz0QgWwjvF2aN5G8
mgS6Pwq0Vz5S2Mp18crHRfATDa3URIS1aMtMsR/B1ceZvtfljUrIFYZ8XHipM3KPizyoHMTW++FS
SCfi+FkPLi4Ntqi8wjvhfWXEDbN9/gKcy57+H4ydh2oPGx0u3ETU/Ggfx45ZRBBNuK+246+/atnW
TtWUjbBNjt+imTfpaDl/9din0gJSRB5G4jSTMq1raFDVuLadgtNVkSl+h5ahfiCR+IdRlwKe2Z+t
ftPKJfQHirnCrRliTRThI5o2Na0JCPWh3Mev9kpAIZEbCkTpIYawu47akqwRyHJFYFKC9/NdhyU1
sYGsRHJ+OqnllVgZ0LjVz2RMxDvdeok376bFAmE4ewA4knwQUopxZSWaAbKi4mRTCMdaPnA4ILWh
kt6oDuL4lKd0BAk5cuDVLqfqID5lhchYcQMwu8nrX2zbYzC5rBoSMSXYkrjk05PmFmyo8uOri4y4
QnCafo8Pq2yrJdInBg2YRifc8kENjJSAmHD3+R0ZZV+Xi1LYkkevuYO3fiOo9GHbxr3zn5eN60GN
eFwxpLkDduFMzHs74RidANfjkJCY67idXxj1ujMkUgU8fB+bYvmXcWO87omLZPFd/guArM3jAtsl
6ah8C/Z4AjFSzuN9NwU0ST5VzPZ0s6yX9ktdKgxeP/1obv1j1ZLAfab09U9AD5dEMdh0h4Mc2tdi
l1e3kCKc7IhMk4rvlwZPEYKpUznnmxYTTgb0t6yyONS+DeuDUKW3xOm0PgmEcFMLezAA6XBiiTcq
UL83RqYMiJ8nNBZJS9fTuBssBsxEsiwJmTfmbBn1TVp+0D7RykHh3cI3uRZNlmcHIj7X5KKbqBRe
XjfOYFIS+z7kosMzv3DN8YaTzXBY8wOD7FKUrVg/VwA2puw6Y0XugA4GOpikwEAb8/xfts0EkiMx
89ik4iECjKZIaiuzxb8z4rDvtGwOZNlHJrjpn1v4+OQbmXSdkVeS+Qe2SgsYdSsupGTg/xLxLbmt
dpXMALi0FBphiyRljg+WIvCIrIGRooSOYA4e5ePudRwTRVwDyqKqznSiuO0VPgn+CSr5AbtxgfFf
uPCC+8Xpa3hsHno5aEuCIceu2PfSR31QO2qkRBH/eqdb3nB/zinsgyeXD9SuDo/LsVcbmYDQwI4E
P9l9aPe4SAddLKX0KkXZnjKrDlbdJ4h9T/NkkigllsVYiz5XAVk6E8OgEGoCVcbYTrH7ZQUJNh9K
80az1Tk3+YJedbsa2Kfs2OYJ55sGfpZEh27QFagzPK/W3Q8w81ANI2xG6DgagbIXZZ26PTBm0EvT
zlU2r0M3+8MPE5eMs2Yc1hVsecMY/3K/htXiWoErjbH7qJuTTcvi/rsiNteGTSmR3POW/gzxDYcT
1R2TzDUBh87NVfaqIoZ1Xe3OVGGnAX1U5toXr8ZlFvmnuFG/eBybqh2yEPeHVJVi0j091t8vI2qU
Oi7QlxgIAx2rmISzXpsXPIReeTJUbaccKHpPSLxtJyoHDiLqRJJLRKhtNrA39xYngcZ8jWxVTVwM
z5NJiXJMnHRy5opuo2S+CCKsUDXrC66bx+qu3IP4juAj5QRh4y9FIXUcjYL7Em53hh1tf3Pobwii
bNgJxyLLWR2DL6NfyMk/4v8scodTWGBVrEINaJLcgpAGWBE5eZUkPRkYVC2XAcknyE4y9FgP166D
NoB5jMXwydaW6eG/5/+jK7cP7E48hP48lJVWd7wbyT3kVdaH8wMYzTiYQeB9HxS3cYzPr6xk5PNQ
MZA+hXHVqjWzWiEkCrvVd6KdFD4pfn+mojcuhL5zrsK5bg0uHRNeWdAwAAm8ABnjp120NauRMuIx
uVLbgiQmc+6tGm0w4v61xWVaPfHJnwyD3DY3CHMrw7qyKzfVCb/JJRKe08cX/o/qPmHyxunuvfCd
MAYKFz6ZoIULAIGplBkWVT+Af9XzoySfbfDIJTRo2sHzAu/YfqSlVR5AOUSqfJs7zkbIYQOEuLTO
AWUWjhkqwcxdRvARhlzf/kj+Bu92LLT+2TBdfOniJWY9HII12wNbSefYT+t1mDmwU4qn6y0IPtYc
fUMxkiRyMJBAUnrkfEyB88453Q1gp6fIDkGC2/zhltfN6ttnALIHUAbu69NiHcLmdLiDEkUzrZIm
tafq7tqpAI/a84JlL3OYyLcVk+45xVQJstdNwzLjtePpmlh1ToaarkcgU+pf2XhI2GtB7wIlnU17
ZQP5fs15kVyf2lGsNvAHbE4dI1kVzxqgncaLS+GtnFutEq4Db0NpHbXz+Vyj8XEHLliFGLlUe0a4
U+ztgZBXVd95ZoLtxeIytokiVCrnMAPrUSb2A7JY/e5xLGKJIq9ijfNbj82tSoNjRKQrjYybMGgq
rEtxTYFNTH5xvHEf/L4+r6Xheq3eOs+tL7RblVH2xjd5QjGvKGGdwpaMxs3WKvmHbUoUvk1tORrK
lPIbwl29MgSy3GSfhIpcSLuRvtD/SYn82ErKzIkByexHFq31F2YGQBIbB60Y3+xrzgsaeaotRkde
upWJUCpES8dHQiQ/ZQe213/PRyfRbCIxmEN2QAu0+CCpT7/NT4AeuCEk1DP3Z6FrGvwEKMxkQMl9
m15TQ7RDpF94nGb5Ab56x02FEX2iHq9NDvlN7kRYSgTsY1YNYB6KgTUZyWvM0xBFLFcdKl1+2C9d
GsSNBPnHqq2mMEY6U49RJAtRzKWaD1WeLv9WYwjLhCtaLelisLSkaspa4ZwhNsFiDaRxcGjGP3oP
VRkcAGjt9gupgCR6uykf2LZ04jqR3TH+T30zxcRHaqL5y7Lukc73e5Q1AgNOd09jP3hopxEfNNZw
5R5YG3fJaM6kOabvx+RbaCsbnH2T10AzudwHqw/vpHt3RFLGa6zxt9vtWUmzKgEfWgoc65aWz7/S
omPYbWzpfGdgjGEBHz3RUTW+qZUFt5n5bKy7sou1HJoVO3bqXa3c1I+MFnIrgMFOgnKg69pBo1oV
00mC5seYwwBcM313KO3bIOiX3cxgXRn4bcdrsLaC2Nd2kqMyBtC3pV8W7gk7pmKThHG4qWWZuk0i
hHZt59QkTEq3ALr7EQabu1boL+czBf5WNBrVZxxkYyLxAuniyBqGXz3FroWN6rQn2AuhT8CP8KpZ
3ftsDUdnLFNvv9GuhCwLIoNtxeZQAqfKsPiCJ5JNq+HvA5kNqZAFKnmRwcC6Opl1EdpY+e/Ess5b
H+5S1ULLo+TSGUeMNO6/Ma6ULBQyVmTEwHZRJMQpM1ghnvAAdp/7eEABsx8ZypyFdafOimlDjBqs
bFO4eCDaVh3lKpUrZmr6NnNSh7uhMs9IqsEIcAbEZwsMIOt49InUdbO66vrEk5wC2A/toB375dKK
Ik3qeSJlYA6H13tlBjbf0Knj+Y1NrMfHN2NBaEEsuqUaRCdw7dee6ov6aEmFSNmFS2twMA6D7xnU
4hSfFykC0kbPW8yq2RHtB5yETIyXcvI1slP7Rwy++BH3/IhM85pzc05i0TxJiK7ZjZKbSxGvIK2h
Vh1mDqsj2vyX9jX1a4uvclcDLh5j+VvgWpXUGd1hvCv8xrVD2Z0BPgs9Gu+/2sgPtO2nYj/nJ6H6
y7ix6MlBG53JeoQYvs07Sm0lQ59YRwzQ+WflFihZ3lyqyqkqEwUzqCpN2ecsr8okf+EMvw14PCHp
pm3nWowsPztT2O/pyUQbb1uSxm855HMPaid7s9R6694j+UUHBlrQPjXX+f35D0qq0XYTMecN79VO
k2CiyPi2984GL6kdkD9OZnWAsOo6LomoY0MEK7baXQk1vn9b6+lbBbWp+Hz22bgWSkXcC04bBjGa
g/k5NTPNd4skgpp+QRdTTYHOe4YJyrlvubdP8bveRtm2uSbZenaaNMmDOoajykXbA305BJyZeqOj
co3SqacgbxYS1yV4ZQm34n8Gx1n2X3MN5Yu3XzvliXSUohnQcvs02dlYzOb5A5VhYfhFOhKgAQ/F
KhsbsnnrzfljiAff/RKHLktB5Ox/gvAaL9amhGbCJw6M+DQt7H8MGb29G7+wBa2DUhERGPwHcFss
ngelNQofJySazSJdeDTu/J1QADfHdAzyCARimPfhXTdYxZRz1mVU0u+i1Wfui7b/uimFZxJCO8D+
yix9UYBkkYrU7Ppq5TW7SR7Wo1xAJAFP/3+Xmt397ynBdwiV9hnixgmZQQ3byGc9Bj2Am3dakvtE
KCoLFcAbCczq12f3rnHXXevUTjAz0h1AqV7LZvTjOAqjPufNJHhqcClblTYB53Gy3ykPdGufbcXp
doQcehjlDqkzvAOl1JS60+AE2USNk+nNAG9RlZ2XlEU/vDllI8entP8uzYCnVPQAs1AIbhUoJvZq
fgiKsBotySxyRcDVDxRHB7cJup9lkZas7ZhpFaA/iNxcRMxhCcqxS5ywGMVOSSwa6eQgKSGDQjSK
Ea9Yb9MEZXKOsBLsGQF2V32j6/vETXByuEZs+zRDzeESPx9AKCICQjnwwJcFWEG0VGRXoXQ0v3MP
mwf+pXP8y2nKkt2CsD9N6k4qP04WD+TDXjo6Ix0gMMH+Bq4LJnvmCr2NIljR/WSlIAI8BrcMbfqY
ZGm71Nn1RoCUQdgBeFgRYeUxKcFIU6O8FQnhvvVMM8iJX08vsoVROTQRPAwOeqMARD6XreyusdHn
8Z/EjH0LsxM4yu9jLfUigMMZ4YsZidxqRuN2fkJWR9mvFzwiN0T62/PfPzAFZCMoqo8E4GjiNenz
SINuWDrnssBta4zQmIYZtPEsfBOvkXcMQED5YixzoONu8UYLsjsdYKDf2ndV/DGsnMUBcR73MJiU
8l5Mues9zFjeo+r/0+Q2fpyMVR6euincC/MpVwYFbQPn4lCQO8dZxWpnZKIq3M23KJzl1mIc07S4
LEqunVkWeE2EYEmLeRVODho43hF2K18ExccvEEz6IdJ/MxBAiEB5nVNU8WHsc0hjRqulOfGtpruw
/dcZq8QSC1JYBbEOIO5MhXYnVIBeKGQ0JUqvC3UKxOl29IhwsoiHgSHwrlC0+NihzcouJRV8nutu
adKip92C2MfzpcKmazjntz3uZ/DsMXtwlwB+vwwmlxNPgseDTjOxNVU7/OfzB9JAjDjYsS7cU3+w
jDihK9N++k4ppzG3b08EbmtU/Euv9Dfjj2+oPzQTdLc0Nbaoh+3RwTjI0JKo15Lt9UP7pk/RYaLA
aKZXhH7tFJ865CrZWwbyLtVgLipH6cr4O11T5pq+G+C81XAOR3Ouq717hVlyXZZRk4Gzv5QKZEfI
nEVqrvBHgc34ghiETjHJvP/JniIZ/KCVygEmpQKfIEVuwoUvxYvt8sRNrn7wKDldRYBYYlACSqe2
R990Tvy1Ha21+hZv0t/q8htPr+DIGkCbgaut1VyfaI1n2Yp1zCEgRIe4E7Gyehs0HzHtoFqRRoVo
WGHWyb9rkVdvgYb9avnRoC1L7h8EhL45+k0wymVrxTtjOfH8818VLWYf24mVXgihdosuJ1Ssw5Sk
iZZ3p67KqAA5xuO3xRM/nXe3dKzbTtYHBXNqV+ssbVSbLYJu1Z2fJw60KrSzx8W43BY/so6wH8np
btCzZQu5553jKK4o20Rd9EPmsiIghuXp4p2wgiKgemjmnZNKpHMwkQvp9KrkkcGlSxaFAk/CIgui
VUqsMxtJGJO8T2MaglYEpta/1qbr0Lci3vHgpuk4aQ3O5Zlx9eM4Du//Ro7yPzOW7R2PiCRZipi7
x005q63h51Sb52G23sOjFB8CG/VP8bGph7HLrJ2VTafQz/rlrjfPMT4W2n+Y1xtVZo7h/1WOVRZj
4DQmOlSSUHHhWi8dMCDtDTCw/Vzl0icNG4RSXS5XQkI3rm99Skj+QtD37O3c6DDsczq8G6erI26K
RP5UOWMFo09lwBiMBEWEDFbr2c4VyU5bmKbqoel+ofjVHNvHagHBVH4CtbZFT6sJZbfjvBUNYJd0
dydcaz6bgEfAbpzduYtsZI2qq4jqJe/GpHl+UWt/VYdO4F6EMapkjA+PVxOOgMdkDoWcTNgltZ8/
/KczcW17xoi4W2KOkvbZb2YzV2sgAMnp0DW0USBlctoS+XGGof6PdxZg9hwwy9SAxL7+c9BbZdTv
780OJw3X1kopbl/frF2yn/snvKMwq43SCpqBMxUyjdenMrzVu9dsurxA0SAGSqm+1jIoh3c+4w0T
D6GDqQgE4VSORFTz2aM/ulFZJj+7UKc3FJfTbPdgZwGFW46SsZU5/ropUO1beh8ajNjZdedoLa2T
Eu+fjxvz67qTDFO0004wCdu7dbrMOB8+VaND2NnSyQIU5vn5Y/DUmbs2+tzxbTSjUjkY1l10+ogn
WCYn0lzEFNqmocDmT+lXBDPPFP3dIJ28aECyPE7YRmFVfkS/yoL3NnI6mwjJWhVkZd8vnDHCowI1
5m6+XVnFgzDMZhl0WOB+/q8eaO/vMHEDYkBmb4ZxGJD15dJinuWYiiHvaEIlExLZegoPsJPr3UNJ
sjuKcckGJH0A6+pw3eP9e4Iq4HTHPBmoho5PErfyqmKEsbiVr1e/rtZUwwHPVERRGAGwgReGtK9L
p1Wh4fzBLVJ7goxfS7XJhI6wwv7LigN+ZOxw4e+ik9NKs2pmZguGf6uE/8cALtyEw+e2BZpLSFJ/
O858VfhOH/loIC4q0PyAqQmav9OIUEuI7B6msengjttvpzoGE6n/YrZKsJvXs5dx3cpDrvhcEypM
aYvi/5i9Z/4UWwI+DfocpKKO32Fon1dnSIun2Xv7hlrdlpz4IbR8lyO5Ov86wSwA6emcgHzV20pD
IyJ7J2bp55Ww++Qfn7qXuhaz+insvg73uH8lD1lsrIYS8kjT7gE6omF6LM9eEDFeWTmpTwRD3i2H
1CHtn08USiGIGRjS8TKfCR3l2lNOHMnS/yGbq+atlNIHBBCwY33COqxjzxk1nqFdsMWxnQen1uoR
K8d1Fn4zwfbhiYNyRtkEb7he17xLYfi3UB8/pMNW9s0jW+cHGD9NIyMMfstIgRIMUYGpYtSFInek
yk0BHbxtd5iYhEAKi86uZ+5YPTn96LE6vemSj6Xn5FG8VGYf//vCMP+SNBbHnCFKIlACbQSUcEtu
uCbXc2BXxJYW30O6wGVGEyXC2NbuweSS7T0UvT2zjIOZjbt8sbBfnDts8I7sBokdbUnTD0GlLg3G
SW8cxwDOmctcX8yP9prG04fgFl33MI5tK3R0lHTGSrCPat/EgnEzvQC6tj+ag5NOXqd9tu+WYCr3
f6/TOpmmhGPH32nKhlE8jVoXFIL9DgCqRAOP0htJJD87Q1QoLZZKvYlzb62mkohEGQFmTx/E5SD1
nI6nXF58aaQ8HismFsH/HaTUULhs6Oi2xb0ghGUGyhXYOnYPEcETsGvb2j01XK62kQTqF8+ijWeP
oBb3vIsUIMKFihdZvrz68mBO0CVaJ6CN5HrxcWPrduNUKjQGse9HFF5F792CON9Zg8Bi5lhzXw7A
O1DmMPHZF9KJqpEXIYsm/voy825rhXiz3ptyI6ejXCNhHxYy1O4Ze1waDloZAQ6eRRXKJjvkOaKr
cOTLdjX12l954LmxqVTc4qEDrKI2GOEJq+837rKooVt68VuQtJsVuQLQveDGbjNbPv3HQ07fqDFr
JLaHPOmK+stxNPv4tIYT0iJj9j5GCoXAlnJhHcSqBbQptjolMSebx4AUV2UOMoG/atVLKvyaCRy5
ezZskXHkjPHLs33GthLaCo2LswpeNLScLnjCeWqU0fgjLGevVtF2EK38EbFoHdm6mi0gAVlC94Wa
wW/JDBw59HsUqrrQkohn9Dn1xIQ4p7XqTkis2ZWCU+2yCHFbR2PNdeZw0wYKjGXqcCA1/HFOt8kE
pSyH9+s8e5Pf4vQO2beHpivKiq97foZj65YCqhoQeZhR59G43AUJa6S8vRJPynl+axFLYbvLle5B
3qq/PfFPCsWODhkLOhWNOm3wOv4GOqejzPRCni3Zm8t9VoupwqVy2r59q1W40DydsS5pXV/8cf3/
pV+PMTkCHFuNVgyAzhR8eBB+eaGtpq+OF84UrOsNctIpckybCLxbJchrdY5tqj8hSkGwIjtIzFn5
wmTxgdCsCOdVheBQ+rCGZ5ntq5Fwbmr9l8Mjs8LedJQ7aR1gvjSt7isvcXFub9UciDeKYnxD+iSp
+Ri40CpQLkNA4K1ba8Vm0kHW/sPgAFrl78G571m9ioNaDIkwkABxX8DsV/rjxViIFZhgWek8zkKu
4KOcpPR6YejByZK3Am09Bt4/4bbLDYdiPv18Dlc99TR1+4iz5hBqPsCUbNxvxTQQ8PITSpWJX79f
cYo+oqfJPRjchKtPLkIRh8jKUaXXcSTOqrEjKssXGC639cAW4n/TJa+hgOHdKWWkmFXll0XOxKe8
sjZo83h0hUID8kRHD7QKiOvkzhxDhpWmNw6slq6WACvrFh4W5Nmki0yOhtpuDGMrYy9aD2vEhYDR
3gtXm3ahqjwHGDWKDVTI4G6Kw869lSUi1/pIAvbpHnIEONBBOkCvF4FKWzgUKImwo8+BflxQUyYR
qBMiq0/cniLaNmjW4NyinRoZvcRtuvagqEoqE1sqmobn96lZE9tqSTHfg4QGHXAYWz6GHxP3RzJD
SQ0EazZeAm8v8amoFuI07ZfmpRJ2QpEWI/Bcw+iRLxiTB4+ZFqBuATGdaEjiCzHgsfkobx+/3MYv
N5oqy7mjJrjokoGH6IGgRHnGLUCd+wi1nX+tQlAtVfJKuAb9y10yua3kkzfIcLROozQuUMYeS7va
RBl9Wz+vaaQJohXLA64VMovYJMqxwbkDWppWvMZ/XB3bOeP+6iSU3eQJUAc0ag91ifNf4kX6LWpD
A9UcCFQwfpLmPqZ3EfB8BkWG8O/3nCFSSr5SamQFi5JvvK6+AK1U5/tEZialGmGDn9slJVgLn1AS
vjDapCGB9yx6Sto0AEtrBJ9A7wLuY2Q0bgG8eT3Vva6ZOrCqTA5eA2/eK6PFIrTBs8zAgrZq0hIr
terU1NtO5z70qxUr2b1hy7x5KW5eex2zbTd7+RPqdXCm+CfFPNvc8/5+sNZx4zMGcxMezC0EY9cF
IgIkV5VpkFKaoq4qT/rRVlb7a7UOobtwRDKYQZIqLeNITUmySSoLQNBle0Fij0IEJ/yasMXf9eO1
pINvzCiRhqw+N3JU4tR83/dnZa+uJ227wErkw3FjpaPov2RJ8Qdgy2R7N8ENzTNR4AgrvJbDt2hz
lnuXNopg7lQGi2aK0c3xvDRA7N9e1u42SqVt+9eLkZVCddTeLNFyKsXuQMJuPU4ZxdkXVP5VdEFq
rEKGz0mThUeW9kao4FsoCQ5nk3l3NhwZRr2weNHf+b2R3usI68F8IVC+ZB+74KJzU4DrsLOlzoOM
NaKusbm3g/FE2W9DGxb17zngO5oOqaSfnAVxz+5pnEohSqMcAgjLDEaW46bfO93OG+HvPdGUX0ym
I8wRryT+AI/359RGSTnmozlU3UZFyE/W8eNxU04JymCY3MDGdtKz1zEWGU+JEXC4ZbkbwfbK+8b8
dMFP6620nLJi5YSFEvFolmfINQ8C30WfLy8S3Cy50hHDHQtE0LUWz8BjlRV7rJ5iNXqky/qrSaRE
7f5+JR2P2+C9qi3MnOtmadmyc8J0dUMAjv01+9VjP6oLm7Ow/W4AWj/lFbrI07FB2Osr8w4e7zUq
RjSstG/mgUmSZ/7Gmz2un7Mv1TZV6zPnBcH8CHIk1G0TUI4MphodE8bDS84Dy8v8H46bQnev+P9B
1A/y/eP83/OsaWdUUc/xoq8LvjzD5JBQho8X1WOWgpTIwTPXkwa5R8Pjfbm5LiSxrAnTcMUJZWfT
tDFGqlY+78/kAWNkjQEd5HoPDADP30z4fS+FYU+U6kaBZxIF4/UYFnlVnfMAp3cwM9fQhZQ8IQCm
F1Z6jOF7lOox/kLqfeSwFHNGwwbc8A+5hHgD3gNrXE5vx+zx7zYdj4yQFV5rDAEPkap1GL67awms
hqxR8W0SGDYiXIapVW5wk8djd3lTlFOWrVWcQ1vrVadfKPEN2s87g0AFgfhu1GqxuSvjoVqOnDo5
axLAm8q6LJGUnXJY/TIpbdPSrJFg/UOFXv/8l3EOZ6U7jSu+dNxXJT1CjwhkA3hok2SMsxqbjEYC
NSugnOIOdzISHCMaJnxQYp1C6VyFGxu8dfb1IfSa55xfuzeQS2sjbX5Lh+Xno/S5mzsyZeJXN8e4
+n5Wj3vdXacV/XnMN9JrfvxV0oRr47YUYE/nxniYxmanM1IrgjreptjvuBGTqfJbaIEhXs8WQqR5
vT/OO6PxKpl6XmNy0vJoG+mUhjEokx8QARr6giXcwNKYgx0OrM55zz0TtBOdG408qY+vp3G+E4qM
EW7yCEozZC3ZYSY2kWoEubAr4b30gG50FO+HgFxNbsbOMoKoQVHqSNG8JuRwxjcePqo76vgQEF3F
VdZxpHQotT//hHbUsGWvsjFH7keBTYWnSR9xjIbgfMtftsqDxfPeQZ6UegUn5ppC9f1FpTtMnXTb
yDkvMKIjrplRROeEZY9YL6+TDObWWBOYzaYriL431rfgQPxsKqj/wAt9SMjFxQto4nmeWXHRh3W8
dQOf5cT6JfM+Go0qgZSf9QHMogJzthmX8zI/a3RjMkEf9m0e5yqOoT1WzI2rXKf+J3uYPd+nnv7U
UMo2rYea0zsTpuJ0EFd8cMQeodWDVtTY61EkaB4uXdkT5kFmYLgSVXCo33iVDIytIHh1OoG5qTl4
ZvaWkEq4yR1trbleop1vD6yW9e6vfDl8RilYSsHMAjdDGqUp6sGAlEbfDbxWIqs043WjcB5I7Y0M
1XNxN3//J4FOM5+x7y0jLbS75s/cgvqK4S2k8XsGvZ4jtVaHn7UonZlNeZKw3QEi11La1oWlVtrx
QMM+3tHj09hjt+mCmaaA+LGd0MLPjv8yJJ430wBiQjUfUNVr5uvjRM8a+BrbomHEbo6zCwQteURm
WT8Y8bkcGj7v9pqh3biDH2I1ACFvJNElXwQdqttzzHGqcCJUnmhgY3Fb+jMhrNy0FcbGnuYBySdv
/q+7nqfzVyOQ3WziWhv/s9EapJ49DPkQNGA1mAQHIOBEAvFt3beO7YxLHvk5YtzsNFisv6Ho3J8N
1h5mrzisdl+ouMWh6DQlhWkXLZxKgEwz+Hkydquu6r6LbxHyXm7OY2OLMV823QcEs31LOTipPDpN
PtftC8xK/1R0J23WflSIpNS8Zq8RGF7ru+vlbwXuxYJxyxDfNdjLLkY7CfGgIpJp6ZP2gZGY/2W+
KkjjhtsydYnRMA4KjSjDwOPc5d7pkctnHP9WH/nZg+Qr8JD3FmP2Tz8UzO7NFMszvlnBpQyudtB/
Aufvv+cYYcbvES1OD4gbLkAwGYZESzGdogmufka7a5bxZ0fG0ImA6joMmmDEzvxFtHRjD1WtqadE
CrUVK0U1tok8iKiCN6dgvL6EtIrPxpSX9Mqm9wxkY0gE7LWeLvzL3TRnuPt6cK1NHJZQ8SoQ5aCR
0oUCbQwk9FPgXFIyAumNuNA4yznA2sKsDkYog+zAh70bFsnXG4xQpsz1A1Obb2ct8vDIU3tcntPh
VmRc0FpNtMpcYNe/8oIokyNnxFH6uF3mw7eyAHhEx/2FulORcHbXq9+XQ8GsmwGzcp9XKekKNyWD
05TNT8lpPnJFCzZ3cNEgBhmwO+1z+/e5/6Houzo3rZecIo4av3hU4hzBx/ulYrxP6NUkcHndXaUE
et3ekNLLy3QAX4Cx0U+Tc7x3a+2Dy/6e991OcGW8XVcxOHIqzGPIctUlKUXVW7J53K9rHRcrIeHz
L+C9rWagwGicCHmdd6N7Uc2MzG+7OeKFRdRtYszDpty/VKdu7ExDYXjSimxzMPBZxmVOl7pi0yvk
hma6WDQvR24IzFv/ASDKfz1okhbkai/bIWqSe2O3OgtO1CB36R8h/RWChAYOZwV2WhD3uVo0g/eW
3vSr7vK/qPYick3WazLh6TBUF2oU7xotr9W43uJii5R4NEE5/K6Tb1Xxc1rQ/LZ6eNt3iDWYsK8b
MxbL2tgCZVFGj9U/pVCcvFllWWIwcDfSIiHMVTFee+I2vqb2CEeSRK4aecnFqaHftlUiZZ/6sb2e
uwVYiq5Wt5BfEf1oInfhEfS1miwdyqUv5j9ticoTZ0ztCPfzFwjDhg7N5kfDZDdyC4X+eMNaGdq7
L/XIJn3XfW0DVYIOE1jr9Wfsc55S7+owMYaI8w/ZfSsE9nYuOoHDCUepgTeuAwKm/VdpNMwPUSiU
VyrwCUJ8gxLe+rUSNn7ugFcYepotPshX1RYTVjJQtASyq48LesqXYRhOcGMaKu7sCGpmSXlotvwa
LjIINg7ToGIBHQFoHfQgcAMWh2h1gAx0/ArmopJxhNqfRY6EftzFdDGJLWV1XJ6lxBNPUA9d1aGx
yz6FpqfKhBPPCTHMQyhqNFJ92Ft/jwnlsXHuOaARW4NaPs8X36z1TMTKwXio2LlskLgsuoLk7Zes
sg6gzZ8Q6dO1SXQyX0RBEQ57sd3ZXtc/4kYoHunuv2H/o+FKblEggOZcwO7UawxxlF38aeYNuoby
JjjEfHnioDubKlm179KFBDGE6SdZxbsGK/UqeI+KKiP6gpQQTnm/y5p/xhZnjCA9L3MxTSk42Xbz
gJF/UasHO3Kl/V7x8gV9qHXrXk3tDR3tGGgcBJ7y8gzNXfrk5f1cQsVhdPHhD/IOvuxpvDPjaBtf
4ZNoCFh6cpYhwpwNt5Zxb04QP9n61g4IId6+4WXkwL6bRU7diYuFYbp+iUZwQWXve2ltOUANM9px
IgT41sE9bqBdh5RscIxElXPF3NomPo1LbslpGfmt6ac+EnidpPQ8W0tbXCmS9ZMO5p79R3fo4QVp
cz1th//XtlaAaI+qtnSFLNr2a/+QA4q1tyG6M/nxGLow6Kj24d6dkarDQRw1eukGnaEoWKKnaAZd
CDrhTxBDbx8w3K/mNIsjYb6sJHszHQfTCTFz75c7ySA7YkQiLodDxr/6tsOmElWym4+kNkrmq0F3
CuzQ4VgBKZmLzHxMT5eP/HYUjZN8YsFy4eJDv9mJXX0mwhTXOQNqOTc/ZetUCYUBBBsfkbsVZLj/
+bo3XMh5dymX0KIj3BLXbF8sPOrXDDfAf5rEKRD55VCCGckqqaRbRg96AkKa5hiytI7MgzbI4X3I
+q+Z6AshUHfEhowoT3kioDT0zXc/LJPHMrXxaDrv3u2FhrwwhvfpGwQc0tp0ecbwJjO7Nk0cO3nY
KX+cYnhObD6Jv0U19T//8wnM8r/yUhd9bWL8GYVgVxokdl96L2p9LVc0UdMeo/2xFO8NnHA/1Y3N
JY1pWPb2IYARrlgCOo0nsGtJYSZU5GxR4WHs9zJegLlQrJsBzT6ravjoDExEykohw3riPvtlTEe8
jqo70ljQC5gSnq9raN/4tqSuBnF3nO5TwoWY14OcBCdm9i/pOOXiKo9V8VcEEBDJn473Ej2l/p5y
2XDtv0DEOktkhmXQ4wEf61Ls3mkVmZcanYnVS9QQdP0U8GsNLZWdnFKOteHQPlt9w/NVYs+Jjxfe
18hlHGBNxftvz/GamFQS6YoqYXLpjQlmLjUBZpGNL2ugsgxYC6IZuOjpakQPQgVwA2p741qZUOAo
oCWpYel5kRdoFN5GOFtCSVUvoIX4DwJ9S+Uzt8ADWik4Q8MgNh1jnp5iwk6nGkhuMUqo4K5WqneY
pusSRnWSbd4QijGWcslqlQ6C5FWcuGvQVpDeJaX0v0c/m2mVNKD0B7tQOAf8llYQF25ELuUQs/h6
G4UR4lgSTDE+/GR31tmEQp0HrC5r9orHyP5lmafbZVMQF3t7YFJiZrejZLhHHlefoYMbzqekLMdp
htM9QW4sKIkpqk+Pk8m8XNvWA1nwe7zQ9Je8EgCnhUfjULyRUbJGlDtRPIFv0nXCrtYCa8Y1kBlF
hKvjAyS+hM3Zvag5wCRsEWvbV1GS5gCIiQ84zhV8aLCaLyZrW0Q7zpsG4SHIRQMp9Y4LgiBtRniy
VDWQindngX3sy9Hks3Ir8bzsOHrzhY5Fs5Fy46gSgr0Aa2+gePcNfp2mVVKdtyQ4HcAX6WQcoOQ9
X+REph0QeBcjXoZv/FhCLXR2oXa+xKjyHot8vw9PL31UDv3jQbiDFg1IT27sNwA9D+JhBU7Lqh2H
37peQlRRdipPshjTaRIiYQ7R6MOQ46OvmAl7/km1mJJJoqb6MGSi4iA+DwtpMLo6ip92ZW4jCfkB
Y2l3FufxuhrsqHJzJiNogG/zPO4KPwxnUOtuWkZO6SrOnjA1IDtKGSz2LvZVoyQGysbOJlM0+ag0
oiSymE2UHJKCIaHPEEmKPB0j1Bb41emAAY9FWMnRxxk55oFbnYnYJJiVWEm0iUUL/agittLh0o9u
Nha2MuTEn1O8VPKo+igTkelZhNgKgfXzl6Vfd/fj+4jcIil112dgRiWSby/okE4WHIwioMaleide
Lm9ilVTsgBlBSJM3hoDDHWajfl4vcblXq5zCDdxT0CWW6xH6pj4ReaEgYbxZ1W/r1EzSM2t3VkFD
W98Vt3SY9L5z1t7yvbM+zHRhlJU+oToSL97yPr5s9KiWv5HB7pmszagG+qiB93j74ExVLwMeXaN2
TlEeAE9ae6+HRGzwnyHf+AQDYHs24uSE4TQQV9QgRrj1aRV3GVpw6i/fj6olXfkLla6Xk4sqMFSE
XLxCdVVVCKzk+65fgGZo4rRyuBjXM1vzsVCELtTgG7s9Svr9AaZWn3aNiB1/RGrm1Vpw7PCGiYOr
IDq8YS3TOw3UnKOOWPaL3tssVhAFDlt2Tvae/rF4UeFFWh2aX/ASxXWgHVPsElnzpuApzEYkY1L9
AlDhl1ejyH77dBci4BiV7n/wYh6Km9gJz3eiw1jRiah9/Od3YNHriBaiDuP0vscMxY2L6/oU2zrK
4ajUvybLF95kupnClbXyrOyCvaWm2ta4aXn7DYKZG5gzDt0vpuRiBEJq8/FX2vY5QFp5dMLpx1DI
vQfDon9dBPOyO3hOiEiFsrbhgbr5suvz5+8ayvq6FV2onC9EB2gi5KILmQAEdLVw9sfna0ssyPcE
AKcXbEAM+seagA+7bifji1czreH8P0grL/2UPdi6NNj8QtgfyteXGb5bl9lOgCO7Ig3Ryj4kDOT7
4dk5RCyQ1bphELFfJeePrGIVEbdzAM00PGy1M1GLXRL/cwEVTvJhBvu8o094zDJU1sof0ywBLmib
A09xpGtvuCQ+SNk3xaFSSiQ3Oj0NsDwDoKjiXm7Fx6K2qV/sj1CXi5kD1+VSvaNflntbOl+s1Ch5
kCydfohUSDA3E7KeAhye/MjK7labcMmIOZjR91rADmydJ+EYSYkyYqR1Jyx6O+DJCQGxEjmPfRw8
pHSDGplMzCco5J8PTUzTlEwn4k5aUee8UTjw9jsp88aP3Anwi4yhHtM8TCmMQv8Qv4FBD1YJnDr6
lE9qkcOozsUoQ+wqJI4PjeGNX4HpzW/gZ6nbGtvNJisLw0AslZq7a6cIpKvEJGz7DDnUM4a1yTYR
rood6JIg2Vj9pmwUkZ5gqVfUfxf6F3rCZJYBQoq6WDdVqjAPw9N3qwklWiQPzC4huzhnDcQW3hYo
4vFGIhOAEX0VxN0sWQ2J59QNKw1c53uhi+3YJGjyKt7bWiB1EIHUXX/hgZC124q9eGpuLqQtDtf4
V6vA+HjpVaEZwV2sURwrTkZ0I2jR6npIRwKuIfrav5M11zCxWxsI+WVi5Jn7lRto18AqI0kN+Pg2
mb/kUy/amwDC1kuh8rE1DsGz24L71M/Hv1kdc2zrTD0b4SgdC0teRzkdt3hfgNH1wFv+nU/nqOEw
RSWWgM0ddXitMYcmg0gTo2o9P/KyvLt7RfpeaHfGlGXIwBpNn0hV+tRHBjAQgK0Z/CaBobhAWuMW
tkAkl8+gOA8dIIGme3DURZbKswxTqltg4eRLyaHDwLxTzXahBDrFOb8xbt8r5CXPlOJX7HbqVqA9
ZIWpGzZ6+amouWtEPdYJ1yRVLTgif8YPFh28Oj9Tbzl3NGiR7oOsS0IOMf6n3vBDPqz+a82fgNh4
zr0yE6IF54IUCjcmuhI6H6XBxJzuG84AGhhP1L5K2pDEUIao7hRTqce6m7yNFGov4pzQrXbx/vhH
zB/ZYIbMIm4uDwfAiHLuXaOvKSgo7cHWZBMrwk0q0+2PSPiW/dJJ53/Xt/93wOiRrqVJF7yO7eih
fzDU3Zt+M8RcmqBdZHpsfkwtI7SHp6afRXkPecSh2IHYrqa8JFqviOmHIX8uXB15FyPF0QevqyPk
9WsBqdtkSEAFP/Zpc/Ewp4bB7vJWBW+oCpKpxHIr01bYKAvdffvLGmBsKJ8ToADFn7Ed1Brxxqi3
uTk9wXdEkChVcYvIptcqP43RX+fMxRWSxRaImN6PehBcnR+dSelGJVc0AZ94PAlYAxdDtI6LPiE3
2dmUDrs+506fNarYjSA74FPED1K72I17ckpBcI9Toz6mw0ImGDIYVgJYq4Hbv3a0+/+7xMyO8pzB
ExQol0qoWQ0nxfcM5cYn9l2WBC/rGBS75iylFvP5vXiLrlO50/IjLmbjJKkN9SS8u6lZATHsAc3X
BQrLHh+pzb0smSmJb8vxFojiVrq0WP1GI2v9uLY2nJj8AF5A+ixjGWN3KB+4+ofZdYlyHk+HtuAs
xnvgVwCzN09R4DmNdMPDdJKRAe1ZO70/KSblWzmiQyUOGdRHSEAdRxiC/9UDxVD9tpDMMwaXuSNA
g8hKGGGNe6mn0d1dzlcYff6i1OtsAbl3HQLIeEuMyX1Y+o6mBvldhQkKis7KJE0E9WHuk590h3Nj
AQJriuVFQDKMCaVa9zn5FsrAeQddr+DYuwqsAHC96l4G8T71VCnTv2tQq4DN/8Qwfgut5tr5K478
wtWDbdtnITBBC2WG6E97+K4YMOi/s9XHYT6GRfZS187HkznwlWShgKcObQuMxsVsoNnfrjfSC+Gj
7MoESAcw5WoM9Yr60O9/xznq3SXy9o1AHrNkdv1x3tpFouaQ6T5vizpxNctlokyuCz1nZr4kMkTj
EUzo2h6+wiSp2CFY7hgRrXhaAMRgiDzoBCtAQVAxYmvy0laZjHp/SHfF054eRUoncbJKKXlPFvhG
1M985pt/E1wB7wbpr83Tpzajzed7BSQbRRuIRbJFKDsn3t084f8urYL2Dj1jigDoYRNCi4Th0mIs
HIm58bsQpisQyQ1a39yHSfHEJxfPDrFM3CBVMO2+gqCmmEmu3T2n6jGDZjKPEnmwL0j9A1/WxpUX
h87J4WvgmkIq5TFwU/G6r2aKjQHKXAMNx10KNrbfmsmjwO0IIXwfwa7beGrsltvK/jD4OARx+Q5D
Kqa2M3biPI4HYVI3lf55nEKy69tljr6iIhKtlFj9rT7ETQxG3w0yloPjXCO8hMVZbHt5+0kkm00A
WEEJbX7+wta/a5IIJ1s8ejSwDEPiTnQxJInWMDTyE1k4h3ihOIjWax/JI8ZZ/L4/ywk4zAddpEMY
2NC51KN7cNW0fRC4fG+V2plKzw38L/C2f57e+KxsNXEBmvACuj7G6ZUB+rbE5h3FDhFA9UqXOYms
yobxdt18ZvtLUdvmydSadtkNfM9XrEfE43ilqN5H5EyTDy65uMKLEkpu3pvSggZOtXqxeC1tqcWc
F456oM7kzlnO0jcNFLXXgSX6hcIpQ4llsPuSw+a+VXhFwTCUsUCHNWqVH8GxvmKyoP3+CYOUif5x
hmR6wo4OTbv0OgpmmE24/Xnz+VGfSgO7L9PoZ8YXtL8T5LCyY4JOQwEpndM/DFptXvaO14Mya9eM
bH/QRYFMY3nYzK4SpW6YcTWP5t23x4VZ1F4R1mBq9GIMlISRAmmj762VsC7iU9kz5zfb3NHT2SSt
ln+iWoaalTjQKKxgjsrdXk6ADskDm0JMKDgWu58eUeHLYmlCcjerSTmAT94fRTQ5JGQ+qW6zkK6q
o0phiIHS0KU8pysuzjfSX4KZYhYTX/p3ijFCftfdZZx/6pL3yI6tARrRR4FW2ec+cmigtCnU9ddm
EtixciHQlJIffhSMz11ES7LGM+Rt5Pq1MTtVplZ4oGWQA1kQISO0+4w8rNH99oHwFuGuvizJ/bF7
7lcN63eClrA1gL9o/+CVLSlXXu5P5RXRz6pQSPca5oSzYqLS6+0i/zTPN+fvveJrJQHaXvWYXCTP
YhinXb3WJE+TOQxBzSfzAEBeiTEpFo3Y+auydL1+Ti33qR/z39kC2vQDotc8u91HBC/W8iHH2ecT
Kig/gol4cIVj7wEGupMZ/DyDe5Rgk6whf/y6q4xUkMM7DeN37V8dMmusf8OoTqLEdPLBiLsb/JDT
20vjbiZ1LaMY83Elng9YqF49rs4WV24xY9yjrsWlzFpGfsDe6kIwxhMcVfEjU0L9Eame2x0FbI7E
eeFFGtyFhljP1Eo++Tpqcpx+cABgp7Hivp6F0rO517o0BDL9I+5Wn5moWdXmwQz0/MK23n+HL2kp
T9VrsBVbkX5EUhCCN2gZq5RA9iXKdlJhj77P6NrZkZGAU7iEInyXgPz9C5k3nfSB8A73S6GtSrAl
VeoByBNAX/tE0RW5urws53uqIs7rFr9KwwG3U28PnIkwAtQPZYqmVbPnjF7PF/5Orbgt00s2lgr2
KZExu2ONX3Tld2sOhExSPX1UswYewymo/RCcZvZtXpzIreDBibfxOWjVIusNt96wp0p1jZW/tY35
6rAajsAXa7SKh2VDF9HzssQGphrfi2G/RBvlCHZJFgx9kLk6gLDcOFyXt0Qpf7yupw6lNYlQzBV5
sjZKZelJv/+IWFSOMyDWOCCsSx2HXZuaTDvNpdZLHMIv0xpotm48haX9Qec+6kwTx95TAlEGdYgk
FxOC6ufog4Isuwd8RZAGgUk1IZGqNf42WFjl5eSE3AA8JFNBkVU7i3pXKe+XRY0xGF/AO8c7C2od
kKbHCYorLHm4yW7q6iSF8NvwNR3nbi49S+bfk1O9f7k5m5xAMtUBfczNojV5rHUrWfmtNJQ7jkRX
7NWZwD0t1EMnj5BXPo2V6W9iiHMsA2w8+pchF1keCpXYqCcQaqmg5F3rClu+lyey1Dc1ti7BX/XC
5UqbIHFnlMMYuQMlXzbZVmmSgLFE2PZjmINvPweBDjqliXHBn/JziAdXqL7AkLBwy6ZaY9yjbRFx
RLxuHC+OT7CNXxScS4+opB1c/M0a6TXUWlJBGFiQuvCUqqtepS3TqFO9OFpJ6doyU9+3TIaswkMl
6wzom+Jh94d/DoMZ3wAogSygOe39GxTBMCY5gGm+fOrG2MJgi87lTQT4N7u17W9TsR8y9+tbZisc
NzbgOFtGfVF2IrXQ3I3+LqOgqSK+kWpCQE7NbwzBMqnKfx72uVRELCKDOgA1AHo1KAiuRtQj4Wll
yf0Js2svh+VJ2KJr0ER71j5QGQxXTZ09rH6weCDzZpGigh3DcwuDHkRLE7K1g7WYRABJvDfsjGT0
2085Jf3dENYC6/NElV/AUuCc8d3MWk6nqo1fHj5smJeLIiXnhdGK5MQ9qoiEiBXKd0z/tq106fwO
lUFNaIF9kExdjiNwCX/uvqmGUcSVRyrvJ5MqEKF5Z3VHdtPXxERtO+yQGKnxlS5EuFsdgO3nrzdH
qH/Dleij65RNuXe/puGohNToL80+8y2+cbpeEMenPpB3GOevJoq5aKhYdLbacMWrg7C/V3KfmctZ
PKP/mKBoEIkhGxrtcw+2UClCJ++PxI9/4kSr6UKADd//ifUwDYGS2HqN64dF3r1oInMCDb5hQTIs
d0zs6rnGfNHINA4W4zn5zE5jqqEaZ6DK5T1yD0m1E0vykt6A/+ywFMOWt+wGxVa/dq837aGwRxLO
ziuADsawFMMq+0/xXvjMe6ZgPgb7k8lxJFdlTMXM/H+N1J/uBNZpSMBGyR318upLw4lk1t9Kalvs
QNvpOg6/aawRyssaOF7MBrbCkneXgeAkMoALdVKd6Xlbs3nNueJDhdKT0l6GlpmUqdrdf5V79QzU
RQn/v5xdz3qVRgjUhwpSrTcIFACLtTk6Kci5eXYVXUgWPfYJ0CKYxCQ1u9Z+0ky9AhB3yxnH759/
cciSfB3mchSzvd62Uk/P6dh2+FUOvXBd2KfYCXt7rqOigZiEtxdzc2wTziRgJ7SXBcR+XwthnZHE
vNLXk5uOPfIa42spWydH38uDH7gl8WeDcbXVXb+2zWtszYGOJ1TJz/o6i3+WDkxXL8i/M7xrF/av
FgNCx+jQUqMHRo3OSCYJowtDwcxNSrMdw0T7OZtl1H75YYE0FBtDhMzZ/YZHz1HKo2yypIE1K/Ga
CFO2og0ykOpzyfK0WAWEy4+zHwXieU/e80jVk6yOeIag3vDZgwMrtMAQ5E2jmmfQ+50/V2DMfC5P
VXAkzUvLPt2PrhLdFzL/LX8PIFouzx0ITye9r29ujg/djFlARhWaYEbl/+2D45QExfo0Cj10Pjmn
VjbSv20TdR5Lgo/+DYY9d6k9ZtBAj3RvJIBsqSXec3D99+PjNF4CNfccyBYT9mngmUCFQ/iqYAf+
PRH8JxLJaheD/yh04/Yh/5sODwgwYodJ2Bq/+uLE/O0PDCYtgzPjpquKbdY3AaNtFwB+qk/Ne6ie
daGqbwt3iFnoC2JMAzYJyaMpTzOAaQ1O3va9+PqHH4S5/YsESUJ+QdNcHTU6yPU1+uiF+qtLsBBP
dLpi4JjlPYGq8VLrYOlNAsf+YtrkDMeauncyEE6JIXWPpqpZDpQrN08bFZVf1N9khysSvUpWBE3b
1PH4F/beadYCQ8IMBWM8zvofQ8Ti3uS4FXDZkmeCb7dPIpLrCuWq08GXKr77oqVYNNqclLhQGW+B
9oPRYyDQ6yGvuW8t0TJkwcS+rIMcMUfnZ2e1gcaiRzTJeXLhJAYFujy6g3jdCdEZtnwx3NeqwFb1
RKq/jGIv9WRE+W7WNjXVRxVGw1AWMGr33Z8qa79sR1gUil+amJo3Fl9oi1+9BElo4qhiOnD6rDw+
H8Kr3HljyvWriZrKIZWX8f7qeMJNXCgZ5yh9uMYIXh2SGsISYM2eEQtSJkbzrCdwOGPprKckOtwl
xwlZpPzi84Kl4d1MS7EsjdAFjR4utdgHIadcjfulLpwZWKWjnJF/YKnqmqKQrENNZgeymP2NsbZi
CUVyi5kBhScNUgDDUk2t08nqF1CkQXtR0b0mpKT8NldWzC8SIKLW4oN0OxBaqZp8I60ijvwE1jSW
xRHO98xxifEoia1a+VAAP5tajYcjcupRS0FSI2yMn31u2HGUuDwJ00j6iAvN4uCnYnNdALWyW9RG
rbT54OWUoh86DkKt0oC75I5w6+fJ76lq7/5qm78LB1wdiz1PWHFwqJq9mIyUbjVF8Go6r0P68t7o
5PW9eAuNMYrl+xczpH3AlIno29aYjZ/BD8BV5d9xC6a/w0RWbCak512S03eQRmlOFdg7+GxWqsZG
ArElObth2ScXjLm63R6lbaVikfGWBKYCvFjJur9Rwr4DqBdqpgKTBRwBMkuRIatHcepNUBX8Kgzn
j6sbaJ3PksBlsOjpFODz953nEuUlICxW1qwRUBiw4ZUDl/LB7aj9OtMF1cx3GwRfNbAcCo7gkzPt
ksdJLy/8BWyXM5NLiD5qF8XNk8ly2t1eZL8/ZQ3USpURKGgfPja7d4L7cLaB/JaoMV80FySCNZx8
vWi35Ms3ihU2xeYr69q9L3MwtQwlP8vd4IyK9kfWuNYrz9n989Xr/1FcHBrvG/+32W9AV5YtiVnN
Cd032EZro5ZSo1yy2WOgUGg5/IWx3gYLaQ/7XOjioUK8eckLkvDrZp7dlcX7asKygnReIlX9eVmx
Svy3Lm4BYknbm4ozAcZfD9DcIaMduHLZFikl/j5in0AMsIi9sItacmk1SNgDcVknvOQo6XQWNhNr
Sbig2uODzu8RjngV66cS1QlqnVc2d7Ug5PCRxO9DVV4tlHq3Cu7MGf9oUNhaD+1ZDNF40Ad0aYp0
L/mtYQ/evHLDEPQ+Inf34Ci08Ieye4GhVQzVjIXXN3L0RipX+eNLb3mFGwlT41Doj5NLKG8tk9lP
euwQjz+wZfqiKcPcZtzhnRg3p0sYpYYLrUzbV/yCMgOmpqaKgi0YC/iZyPUVmB1oiiiTTmsAxfOP
ZFjWPecqqpi854L/3cKmMjpET6vdRGSgt331PG+oy60SP5RP92oyRS2xUugfvI9yH4xUAYOXAVMW
YAYyUyQRwF0ZMjJ4WsC9a8RY66JzCFxEHCL6Gpxd+Ue0h8gD1JmhN3dPUG67izvnP7jKVVrrG8Tv
QIlkoW4RcArDWvrQIeMtaTn5MQoyfEoghAfW7AQB8n4Zp4ygS9XKXx4V2kklWKZDn/qJ0MD8mpd8
+D/U2v+tA5mESAxOcHSk9ABHptuLvyxZmYfVizjjQmZbYBCNQ867lqLPnyY7Cvea/kFnkATbusyV
O+pVVZcA8YklD07sdsnH1X1uT5il2EF5m+px2mf1b2p3CWktgFqm7JWryqY72ueOAvHTHS/ZCKUj
eZSb2JkP/ZKifGNhr4K2oLCBU3tKrA9fZRBbnmdtGAxVv8TgRAM/r4StYEhB3P40chtu0bB66ISr
nmfcG3jfDUinR8rhQvq6mhUgpAjhV3gTwBQ3pe4/RHGn97dAzeRojIALa//qlqdU3VMlo6RuKEjK
Ny+oKLCrRhZ3Fxh6emrh6B7LpjIZenrzv1qVvH2OTrrHTplLgrnAHzbsoZbHMQqIsB81xDqI0nUK
VOT3KORzyCsrtGZ3v4Kf2EUoaA50J7WQ8W8OUahr0kv7kixeK+2DGnnTAoeJ0PEdp3iWFtbGegA/
5R5HfVH8W96Sap9S1flsYmvfb4Mg+8YG9lxyoGBrM8MTy62sY/Z3upkX0aF3vKzrzUCfJQ8faM/c
rv1/buii0DlfmUD2NqYBzXb7qa5TFaRsvFmwDGBibwQcN9PdJvL5Af2FOM0302KWGcGLy+OGXcEI
k4EKSnNb7+54xRsky0Vu1B5pb7i/HkBbhkV7X9zMaYKArNZ94GNrsPvhMhlbDkrDex1+gtw0a3GG
tCFYt0SHIqEkcX3va8KKDtz3owwurUJYsDdcDk5+8iHp07kFVcz3PljkhPZ7kUhTbfn0TjDMNxas
3tZxuODcLMiMTF3oSpISb4Vg0q+OwO1eylvPPNw0FoB26rZ7UYwd2f5xfcbx8KTbi/lchw7LkCmc
cxZ4KZ8pAZWQDR4wTdRPWp+s2T16Vbz37Bluk+VvGxR51OQPISTEDBGllT2PqLw2R/dWOxOBIfrw
MTcNw3c6Qx4wA0MfQBcGEKG/EugD0FSGFMOcsvtT1GtTC2YYG180Y0fF+lwXntIP0e6beDAiVIyI
oogK6g4vlab2i6v8OeAWuQ5kVrHOqiwHD6Augz0qo3dB1KyFHV08ZwVV0mCIhT5mV71zZq0/Iekx
/EZrUW8VYgWCZ5QOcY8ynxcioq+KpoRLge8QUmVUIKZpxOF7fzlkWvkHC9cQgXrRH5fZjIiFZ8QN
U5LV2jcRZia713gIi1wpvnxz80lzfTdoVafwp7yyajQMmsWlxo7V3v6PpZCXUfN2bNkiQ0e4+bra
4W//oqK0BjC3BwSD8F9aHbdaN/XzwkrDH3mIzol1VYaXebcvmneCfqgkaE5qNmbqP4fB/xyBVK9n
LqU3+d7/Iw8FcJsLSY5PPK+yNOjdjjHcKlIfTMPL2V2rj2Cpl0XaOfzdiWe1d3JRNPu9vM6RqXbO
Xhwx2wNL43+utS5rnGYmDsuUgt9VMo0cwI+PZfuemr8ZV5i2LacpXBsyqkS6e/uB/X/OE6AaN4w0
8ehouTgVlWP6jzY9xwmVKsCwunJ8IdjlEvZNIIzWTX1p0xah2vGXIcUX6d2+9FGQYpRfWBxj5Ngy
AiCz0ieFBzqftAVivyBGr+UXsYm9xeUmB+CaeSfQLGE0LWgUMqLqXm/Ey5yVxPpqTYbhlpd22GCB
tIJMmkzYw6YiRxtQF02gOkjMT5xmAueZ/oaV3Lcu+mNuvGVZwQtlvEHILUTrz/fuTUcClau2u3s/
RH/jLJwxwe3ozIi8Ob3zK1+6Hqpmyr7/asXvd5WFEWJLMiQCKM8oriXAQi3lFJBEjg2lnDRgUh97
nnI/iI2ukPIW8fCCrxtB956WCCn2kf8R1YnlJ4KRJvQaV4q4z5vmCzjPr1B9Oz4w9/3un2Vy7Yzk
3AtPvQl8iDr6XGvQexRY9IRPg8L+kRaBECeY0gl1eNQ1hlc/HpcAAnBniihzempJLO4eJI9MLpMd
nmeW/cFqOq3ZwbrpsCMEzbAR34dP+ndWAs8lQkPg+TmIIXCgZ7o62m30+kR3oMnPFEkAKlDD19Dx
4pWAEBQXD3MHpJfJuAM63YA0HOJVQAVJZVC9R5t+uAQZQUFGlQAnmOONDglEx1uARgZ7H7RyA/hb
faYnyUQrhKVBZFINRkAZAKXtIJD5bqLOw2o5BvlIF2j8+gISNUhMFYchZYM6SlRQlbN5Hvr3/bvG
/iKlq8/n1kYI8jvkmJ4JcvgAYC6TSaNejlBkeF8QQm4pmbpOVadwQOo3rNzecnH/is8tjCbtfWgG
yEaw51rybSncGeKID32wVSodFBo9/+ssKIVP2ZJn6SjqulEHWkWKAwzqTwKS2J5rL2ZJzduVhNMT
iC4IyZE0LhzrBxPlnf3JXCqY8mmJc4y39ua2cjZZ74N1V9JzApzIin/E/Tv76STdxFapvEqqWjdu
ED7x0g0Tc4E9zpOmCdmSL84jUIF8koOw6HJlOT81jdS6/xJz3gye3gfEF0EZBQOZloH5O4r+0PT0
z69hSrISmi+eu1HYqaxQMLR6NzbpAP/+treE4qRS4ur0AmnvMJD4kq0JVzV+wYtE9Gpm3jCli98j
yvW7Te3lLDsKJg4662EYfdWaU9iYq1bXy4jz6lnCz4ELRzNtpr5PoOKQ76BwUsynvfPSqoAC69K2
WCbeD3DRhme0fqnKBVRNU2h2nJfMhL1ojm2o26JKOmsgl3Nv9/8pBzHR6ziCSAPXfuQxux+0R+MD
tpRUYJMTV99MokI2JR8uUHtxpurUXaV0197ypA4KLyG63jwlJlb8MZCPUN2+/WuhY+Nd15LXBJkv
3yKC+Bhd1XY+qRq2QhfJwv2vVXJZUMfUq9L6LblKg1Ejl7taI3WRaxPde+7Z3cu7TCICfqWcy1tp
2KPbAos/oeYe2NePY3Kb4AElJ2JkXZgWuS/5ZkvFaBINJONBxXOSd2tkrAcKeDOtsUo/PfAcVu+S
AXEUUV7MFkO/i4nnyQI+Q0cGZ0GhRDqkV082j9PpqciH0Yc6ntx3kDEnkGUXuZk0LQEhAJz3aGMG
CGDnGz3CI71/Sl28PYvJsY7UnJAdqeloCjXd4UHNAeBIAQOvUNNT4QJAqVVdoGXvLimP1yYOJumy
x0LKYDrGN9giHQhYlvF1xi+oRaZpu+CQtJfV2f2Gk5YZ1eS9ccQ2WeH44gEd8T5Ag/weMuLJtwe5
GeTYNeP2uBGqv438m1N24u1k12Pbzt2XvIAbaJ4ECARHRhVsG+lDcXA4GGaT4NSaTdY00lBRReuX
NunxiBOBVwFK28UgmAey25d66UjrTAkjUd6fbesRSRcDOrU/UZZV7nfIFoLPuGkopB01aWEQWUkv
+S9BbiqV1UlFruqQzXLko/fTFI3iz15ikbtIZ4/9BU72dUaL3OqKVFoVKQVpoYpQiZ+YyTSqk/O2
WFApV4IvO0T7LlZu+TFRCBy3mgpxBa6mw94jMvNaGRkPlBPIOjS5Fommzlh+JFEWYWjFLEXiIjdX
Qu4f8aC01UrenCaBo1tB1fSyg3eQoEd8aGxsOXv8bO0doDN3lsSemv0sOf8ov0WwdxcbCsPZHOp8
r2Ix91ByZKu6AywxPdS9fuEY3Lgx/je/5NsXdN3p9TxZwQ2mWsRT8FaaiwZvLOyi3xM0BNPuP7PJ
dK8nn8gGRh+/JX+X83Cb3sTvmlsc3quMjzBPF3jv9Wm6prL2KXsXzYJne0HkAbRZyrDr3Ialws3d
HS0hMrbw1Fr1kkDmEHh2Eoh8KBfRCiWtVCPfBfJGHZKOAfyX16/YR5DdgY45Q2Ta78ki5y/ueHqu
er4cMPkbIEaCugbP8io0+DzZ0S08jT5fGJ3Icci+0xhNPPCFcZ2wq3z8TLYXKHMc+E4tFzryHxRG
f1EoGN86k74gOnG+dx/qHPZet80bBN7A7uz3hVN2jDNVwPJIrtEtEKyu1nKXDuKIGv6yEaXzAI9J
5UqqD7SzlJZuGAwaVZdPbAa3ldDH5vLAaGc/wal7FfrR7zaLhDqC5VMlOVNeCaBgaE0Y99mH/TzU
hd/A9Bxpqwf00XfdO/OIBa6MEQJdAlpRY7DM1QaqdeVVAE1gn2MVpcEQm+L/cmE518FnSrN5X7de
zKpzITEYS2E6dIdUwigCXwANy+1oQIH6g/wvVHfnCE+LeMnBEAt5vqPj7/qW9JjhUJb6CMUCF850
nhgmDQb5Jzcl698JWnfhgN//cBBkFr8gvMjjQ3bhPU/obbzycvS/2RgdX+kXNGSAHnxzN7OeDnIC
BSrEUFC23/cgRxuPSG0nfnFwCotla0Z6Zusi6DxG45YhtrQvbwC8KtyDvNkmzYziXvvM7VkSyxml
C3mrArM/V4bzcnGTBJbpr86Wgl2kky4xBNL09n9TzAmMTIFKz5+p6cExCfQ6PZwIyJfD4BzO2Zat
SqP2WqpqYH3oWj4zVkOE+cTTE6UYvNd2jcVgW/XJsMEQPc5rKZGbCTroPe03QXufdcN2y4NbaXOL
dvKLEUCzSkE+deKgB9WRKolDdb+34Dz30ZZ9Vn8mWTwuIoqt0/jXLCVQgxScKHA2dyxXuu8zAejq
Kd6SdOaUIIhaNT8IVsY0gYD0wbL57k7XKoN1fIi4CWjy2r84or88MOsLlsbl2vpGE3uIpVl8YOCE
ReL2JIzDTXdynvvxO0AliqX5pCpqLRg66DKpmtQSpMp3o5NVXHzI1iUrj4AEpojSfqSwtnf2Hixw
AYa7JbcYKThvwH2cUj0MBtXeFwR6z+SuMqRbIATSiyOZY/RR1WJYByJqZqOcBWOVuM9cY5+5FIiy
NvzEOovb2m7Ee2ZYY0dsHCWdi09xkpALzNr93LsImCkazPZKQu5o31luFQu3JEXxnwmIIdR8bOKK
1soZwBeHaxzoWThkKf5V7qzX35NR1Mq74VG8GDu7B3zuQCLHxhY7OuwGHFPal7DMnLgpG2XQwp5m
xIR84xcAeXT32xGIhozHBSZNU0oPwDRo+3zAwCrPXs8tf0XAbpBUqIBBcMty7ep6r/0TuW7b3Ojo
eEm7s7+HYxUJsr8YLPUvR7OA0cMRZembakYetUlJ6CuZkjRN+2XEG6Kb0qDpNWMplssubz81KIdK
qNQQ21JK2bbGpYHoVSUc00dBMyyzdTgZmQLFwLxh7HphP27+T+RbHR6l4XSn8WaQMMDLApQySl2R
XThNwXlkPJrfiyvZX26WKVlCo1mGWjttkcvLXcjpFhpo8AnG/aaxeJ3JFXpQX1Ng+tElqXKgA6BW
Y988unIn+ekKpNsDnAjAPj9h1vvglLjdRwh/IyRsARaIjgqiXTVzZgp414rgWs/FaDcrZ6YnDr/s
/NM8ui77iPoZtZHakdiB+jGct9MgW+oxnckTD4xHUI/7Wkzyvx40duF7iZKBghzaFzE08THb2v1p
f/3IH3S4TJwmWDUoE/6MtSAeoJvCUAXvwWos+te0gQWaxcmjQE57aJ5Cc11yMPOA9qcvWcaq7ove
hqxUMAyxT05oPTfswxqZyQckq7Fqzhxhy0IekUO89IvpXlN23JYeT7NTWg0rbstzQdbpoi8N0aPH
HpwCLxRF0pZe4myS/p7IfJ0E5/99Lo1sGlY5oYJvADDOzwCcmMoAiLnPI3ADL8sZdSU83IClDNYe
VwSdk7jReKAtjIoNyVN8xnPcfOd2CeD/nodgR9drgcQE0cqpEQnpb1rVGItkSyrh4cvZpB1NV4AM
bGldXjNf4vJzMchsF0n1MZYdy0mbW7RY3yCC63DxkdO3kEdzboQGEGg8k70veqgZN42i2d+p+mtn
W0HlCiYb+UoihXtAUydytwxeNcZUqCg7cQwgrkQt4YSzq0sEbRbdZm2dQR12eSvtWwkyuYkCCkLJ
Rv3FMHXlD0zbCTMiq/kLNtiDyj5UXUbWl4xnsufgzXkd7jvjn68GTANIEp+8ZsrATAtVrefP0i3H
v/k1MIchBS01bFFZxjX+kgypdo/W6YtWGhurI3OIti1g9WU5Vg4Nu17YfT9tv9kAb6fwHtAWNk29
ybFbbkDnCOwrv6sQuJPBvyF/kxTa2lHYPba8zg009IpqLUHng9gXpKTyQws4EgUT8Ex65t8rwdGn
di/124qfRNsboXFUCoQaez//XMQIFmnULbucJRM0aGcSXOs3ra3GYig9ER7nEMmSIehELbQW1uEY
QfNQoSSYevd7pa1iNVPJEw/UZyQGHikv0TmHsPe3z/6yEilXXKobz1k8aAuya9cn/brJ9QMdEeY7
1qMbEAb12skCE3+o9AbfirRumjW1eUGKHZxysM68ZZpQoBh/YDFghj3y9U7AD+bUd4zLeqnUUsJA
sJyZ5h4/arz3U173vrLEOoVbSApMtRGY3GNClNbtKAn8/5M0YB8DGNr6tr16FMjKC7P4VUsDdMOv
AZU4Sls0Fyj7B6Z3Tg7ARCckE4K2qZQAhuAJt+ttAvAKnRo1lBNTVSr937WP5nq7+YRS6aPpj5y+
hXJLtF7LlYKPFCHparJlla23Q7fQ6Ef0y51T5U4WwsXlZhJb2wyt3y/NLcka1a1CaLaS3sqCZMF5
Rvx6J243eXlMKCUNERnFu9+E0Cy6hhq65qNgAQMhJV+fhtNw81TiOfM6ymICTJ5hM+GTO+ozjeHC
NgWd3E1C+ZmTE+PrdnHI09uMFIUdaKMDo6lz5wtO2+zm6l1VjlgpZYUqbzDEcYduREZlFCFDZcRB
aFfxQafoo3fagllPxG9NF+RfzPTEo+pegtbpA3Mv9ewFX5ielI3H5bsjXWW685nGTgJjVfCM2JIQ
lsJWdsqhIdo6BRdkMRSAxatsPCGUqbkX2qVHyEnXQHx5+Xle40JFnCna3VwCkNo2euZrToJUU3GS
ek99ho/r2yNtF9uc1JILYwMcAdJdyEFUk0780kenHJH+eD5bMnljLRgpXSdhM00M9NiT1wAwK8i2
0KVboGdGj5FIKbEimFclSx1hBJbzibaTOFmsbrQwYjCpk50L1nJVaC/BVb57yX+MTJX/gRa6OLnU
zNDxLwFNDcj2TpGJTqR9JOgoHu3bBHLOsDDBZRExqnsVyrXwyC8G1F1tBxE6EgU34tiNcVkYZR32
dx0Utu+8MPD6/m9c4nJ/uCrw9z4CWE3jmW6ygZeiHBwAi6tapLlZ/lBHDOom+iLbtw57YgfqAxPn
2qLW0/cecU6xK0HyrLeXHGplrf7wYBnZEwn+OqcXhu+H/i6K+vUkUtHTYi/CI/m4wsY64Wwd0Liz
GEEGAOflKAxzDWHbQ1WVUOB5O2kxeiwdpc/nz66KlQRB5KPbEq/ROsYMidng2/Br59cpOISvohzh
YYUYfeqM5t6UJBbJiuY1yAiAIO/xydEKSI9j3G2GEzdgZDTzIcFqNyzCORgVMvJEr9d2w8ZPZ36k
VmN3sxlv7pB9XJVnYslOAA5k4ar9UEkhXKYpxWkxlXsVR8Tl+hYlJF3g1IqTu1rhbUcMTmeZsQR5
Wd8Lb7AC+CXi1Kudp6kP6GG0zyDsty78NUgaJt+E8nzCq/BFxAua9XmUwhFm/G6RxupRkIouAa6W
jxZxu5OewBoNIsfNotgUHz8kCNSxUDTqT7BefpARsXSVG5k1swnBEqETfTSqvzxdXXtCGBX1oPwf
YKu7o4MFp+ueNjsZ1PZEF2FZElNi3q6PAi9SCOppRrA744/phcXzFWQwO+jat/XrvBXlwuxG8IZd
dR151Y4ZpynYi2+AfPPXpVr8wGEZgEbZzA+OnPcnA5XK4469h1Ulaw86GgwBTYTS/myBD0SLMP3P
Qcfq5U5WADTJZvB3pF0fYZ1M1tJOYs7cfs0hehmypJOgLCmQZcIukkb6SzkSvOxUnTlUqKFqGTjD
qDglxpaLWMQesnDfjcWspa8liPPRfoOu1cmGnHTf9FK6+kubvO0Jdl5mfJFN5NJo2KdicoWmif7/
555jqfIP++oTkjmG0OkLrdzxiU5JFMgRish5TyDtNE5lzLiGweuoriS5VBl2u1aB15WqMjvLs1Iv
3ETCkBlqsIFy6EUWiKT7PWbAaKa4hSquf7EHqsX+AcW+1RVIB1rVRHcHwRQN1fPTLdbSvg6P2Ceb
+colM9oFY9RHGxGIZWKg9rpsjQxIsg37dwYKoTl0le0CeWqqZh/D/BuA/UO0B7IwI3T/04nNuk+7
3/312990tHm8uVSMKpwYWHGYkderqVnTBJc+9/Ta9GDDZ7g8KNogl2uMPX8vhoq2Id1lmi31dkpN
jdPOItWmkpmORUFyuY3XICOe7N8qod9MlEJBTwt5Tti2z7XckbM4qVhV99ZHn6rOuoaXLDob+0w0
vPlB0RcpRWzSWpn81qa9Ep+8ddKgpEkbZgZ2W+oY6kqHxY0rBreUWwQ2IJ1UdYPv39SJcOsQW7O5
vhnPVNwhGX5LM3OPY9B4e2wsb7jrHsp9nUAts7O+x5do2n/s7PtD1zRT2+iZUrii7ypmub1L9vNZ
lwUkiW6XqeipJEh2B0x8OVu7hQqNFTiBwbrkm9yvRDej89ACjInNXc/OfzvmaQaDs/BagJm/rEtK
axJSN5LYzn7PuryKHd8oU7cDDaGjE+n2ZKrWzXLmAVvQ0cXjqAPiRe4u4Oj7UeorK4Nc4MmU7nK8
TzTUMCTojGMwnXlxyYq4RFUl+7/qOkfcWEQISwaNn1U1+Fxn5TUwvPC0Y4cvgV4Oo69NzvbMtOwj
kAgmi4yKD59WB5O6e0NwfnMRylYPEvz/7apqTfsUNyPoASjrxbOFAT0dFSw3zXkfRtDfTOmK4wiZ
ruEsEfu5aXcMnrwzCDAOKFW6jjTZYeKD2Umez01LXsRovH25d/T0PMFc/1OQKIs86n0hk0sKAn2a
N/M7z9lBgosJSVthb3d3j8a8/2dbZJ0Tyhlg9/ULMsqw31G9SGpxMW18CgFCOrLe7bxO13fYBy0v
stzq5o6VZ/jEgGmWNiYwZoR75hJRcSse4VcDVd3/ZfeyalmUeWHkRAIG8ynwYWu57uOWv01hJDvF
ppZR8Q5YzEefEfOgDUa8WQFNYeDuydIDh35XrDeBRBa1r1H6yYVjISMuYfOWnaLWj+0YkRNj16hB
MRkkNfxvjPw/FD5uXH6Vkz0N+H+EuArBdvnf+pguTfuEFqFF/w1cVub2AyCWPXKnjl+WqK+j3Hs1
EkAhO5Ep5Q7XfHLuwdOG5AqCaOgJKVmN36EeuXRG76hzDoNcXqxEt1a0XLTLwJmzRJQm+USzAsl+
C0Z5dkDBJI7Ood7xz8btuJTw646fiPWxr9LluHw+Y1wUUqwXbWIIu9ZcY7B8eTSPEp+urkyOYKXb
rzWmLy4SJAgaHmtQXHVjZDyNrw3P2bK16gaTav7Nku3Oisz8HJAK0NsSnT06qja+cbUoScubNqNz
szg5rtr1T7Q7su7scljs4evDQjioIODd6XRxUahlesuJ3MoNYMKWlqYexUbqYqb1P2GeaN+mWLC4
eg6oOOuO4TMNKIIM1ROu7mRwFgE5VkRz/H2jScpCGvDMQGuQX+1Grx6Lc175qDJW6q4IkOYtFTgd
AUMKhyu8mFZ2ArmPO5GTnksTHfLVXp6O5/NZl6xujYr8iWkQ6iOUtvofDjTmz6ww6kwcUT5sxieS
l+3GFss6gdIyABsaGT3E0DARwd81rORYu4WxRg5uLEK2NyiEd5UfNliA5Ao44KRrpW6YpwqIEhSb
HF2+roHx0yyCj774V+OMeFY3oOdKn/L9hAhal/xn0eWOyFp+kLII8BHDYOO+6hKtxYmLUL9N7Coj
3tQZLZ4fkc3UTdpng2aXZlfEe89fcfrIKsiTRy+0XzU+HqSY8nj62xdBCEVEJ+6QNjPOEQ451yuh
oyDaXh3K0UkTs8wT8CAUX8c9LTYOx7S1Gk1s5CNScvxvbqlZ+RgO2bR0ig9a7cpuAXWqI5slai+M
Qjry+DCKVdhJx2UzVZe4r7ZQ3ae74EwDCF4mSmiJG/EA5JpyDQ/TabTK7Mvty36jrHusBhYSSSh9
JqUv90+hrGDBJqOO2u2g/DWvR11kG5uZ7F071WZsA3qh7Xa+QQieKYC5audFEetuUSgmqvhj07pk
tNF+z5lnQ7a/aLIhJBMRE37Fb0zi/CkoqmvmeD0ACdd+DPsFKy6aikxHRKwm6yowRHsM+SMyHmhC
c9Va3FOx1HRjn8tg+VakAQhkLQUyZZ54H98as7q3gFsMn1+n+V7a8Y9Ih2FKyoPTrGCXT72id5bZ
BwcjaUSluOPNF0jdWOs3FfvHCJoUv7jekhThBWrJxmTdSPVTMTzDXzy3gdoKmoyJEZF8nCxESPFU
+qvWwqux5j8O5S3mtt+e1iBE7xEsicsbBCPrZmVCC49MDLksVsV+yXm92N+aCC1+8rP/GnZg44CU
9e1fVblxmrvlbVzlaeBSVAWQkmVVQC6xK9q0s+e3jZmcZvRDvN5AlOqvjR1ojwzBJRLsbXgMvHqM
vF6sOKEqChJ/qZ6TSy76Yyc2bCkbDFV6CWAzklKYYfXYzI387bAGw72erkAQOhSXJTUTxE6S64gv
cEZ8B+sU2U93Rxop6wWsss+GUVSC5F7FXx9DLhAlPK0W7GJfQQp8Sam7FuA0fyfOKQ4+1Lq4pFxY
DNuM2ld67A0LvH0OTUlGvjRWCTZPuOZLxaKqt6Xivl9las/P0YQcDGc1onrq33mkjutKtwDIrark
ZlZjONbXPCdpc7JCyrh04Eff49Dm2JQpPY1Bb9370n5uNXeUdVy/cEvcmgPs+J7+CExsFf+UgB+b
RcjDKwSkyGmqI7y2W/rJ9yefP6sAGrAAiFQCBm1FNmNzKWLoNk0H8MxEwcnIjZ5XqoP2FDL8yDt2
MmpoNOWZowIV3/v4L7O42afXerKuWyEQm3G5Gm8FPqmkrMi6l9i2wM3u/2ayAWR4Xch2txuQDZi8
yLlniiP7UFKYAPnkDD0TsvA32D9pKvvHFOtfXKhvknNTxphe+t6Adbj7PXZa44913XEb0It349pm
h2Qh4ak+WCVonly1BRcXHbkxEJ2sby7SPWSD/yk77uCUz1Ox1YEDlANUeflQzEtmjcwDcV9wXVRo
OcdE0H2GW+JfeioL4qViPcpYRIAmg8EJC9oz5Be1SpebhwNJSjbE605tRpAXiiSHfFjeWAQU37Yw
vWfd5RAJ9udv/EB+SpWIShUDK+WJtA6LCXDr9UcTOA2hqKeZuD9NJJHKRq5OEGfO7/2r69jhA5s5
cf1tIt/0bMoE5EEfvHQWoiYqcTMDOTbsSOrJc6tsRTvPO+rbl68ZS2YQHv7IKqpLdV061ekIkDic
Oy0erDD2MzrsBEKfGDfBpIrWHCn7k7qzbxpUn5FMWe64Fxcl+hTuPgCKjypy5CsfxfPqiOycAm3r
ervLw6L2MVoeTG8Z8pC8U62x55SIsYUDTUUeNrcbgwDzfChtIUZqkc7zGSiT03FrM+e1vopW8AAS
Ocj44pPgOa889eAf4BnOGRgO9q8poRyKAheY587QR5F5hoTDC2Aq+uU1M5nMWZFhCX+8qba2KD+L
zRU2SmXEANBFlSayk3WmWXOKQyXtnjQS8DSkfiNcxhaBTOXdL2TH6vnS4KzDwHl50EJIh05mwtxr
nEhFNelY3AT6Ofqv8WvZnhBZnyRowra/U0rCjYtzlAI4DeWnyTq/7kKlK7kKjZF5oahVZ9/zkAw9
0TSkwNl3iN4NcGWHQpJCLhC/hSrOgBcpI31PbZVxzOhMwo6PioOJgAgGUfjZgREbMV1rkCpwvIar
W2BCI+Ppp6QkfGJVJreMEVCBAQebxU2f3JEyWjof6jKYpYzLSaEEGkDJowHoEqzuNXIovdcwNOdp
hkbqVmlor0VGGCcOpjeur3sYe/fWGW/xL504Iwln8lZ39yKvmcxpQQgYfSHnBQmP229e6zi2SuGk
HO6B35bme/OgzyzA+3AJ05ZL4ADkU07Il1ReAvK/RN3TCEEjJR/QrjmdlUT3Vl/9Tuch7i770x7P
bxbypt3RjKvODJmpFRYbJ+KsiYS7iOzBPi8pGg8yDgvvyHzQ+RMdJyVtHfDlNYuJ1QIDh2oN0b0a
1ZQuzwhClK24hkLMcQtUEnIY4OpWfzDJfzt0cRgpo59AMBULHL66t5XIl4b9wxYVGIbbiTudVFO6
EqOXaomKeX2EVlB6ljm/Lsv5xJQPaJIAr9CMkuEbAxT3jwdHD2uvYp//faRuerd9KnzCKOSFj53w
VARwM/aG/eDcRxD0iG1doMLzee93tsrYzdBdPhTxrXAKDsTOflAYNnxrGAFeAT45oo2mxr+3Oe4H
u3MH0S2e0ICBhKTABKESRuPyGo3U6tGQZT2mlrXv/Nk1mPSQMrlxiui5fK5rbeBgF27MoMYm+Y5p
WOzoWoS3TkuTApBaAY2huNFRwLEOSEHf4dQnS2BW7GCbb4ExHJJWv0zh4GITE7Y4HtoD1Or6Um8/
q9ld+FuWO34q9b6BNDdcJIxUVgkkexWpxU+YLgHOZWZqY2hhsUsT8BR/nZPZM8kgRyJdvxKJ8TT6
Q3QkQcN83KOqNW0Gom6Ds/+medlKblrCXY33wsXEHmAl+9/8cWuZSV9P82RdBOfHjG54iLybJxmK
Kt/EPCxgdkgRiwKmLo9dYsO0OU8wKZE7IXF1lwvbasNUpVPyOSkJfLVnL0XDbsRVCth8iNkdTmSI
FyqnVQIHCSl3BYekwH1p4Ag++pL09UJUYrnXUxECPGY6liXZyZSKU59sdcBoS2v84XwsJ4RFQ33g
kQw6hAO0NPZoEkEv8UNWEl/iywvjLl8k5AQdxhdiyUSZZgcpkhEiTSig6Nnt5f7g4Aypn+FV4uJj
3GuckKmswYKnj5NaexPMpd+DPmhL29kl8keJ+3z/cFjtHJQ30MLhQE5oiwdcwq047ItmPPyF6nqU
80NU4+e80f8sfUlKtsDQoDwPh4y5NngDrXZ3z9fX0ofA1+xrAEhKURnJ3QnOV0v7OpxDoFan21H4
BTFOYUA58RkuBnTC69m4vfpzbArVZYUKd2pRn6BrezgEaDJCe/j9UF1FLqD5xl+GGTLY/pnUZsL6
WiZB18y60QRpCFkqDkUKzUcqDLxlWF7v9c6F4cYTbQf3jUfawnd9sgL2wSSy3zRVfVtrVZ3z5XAK
BudoUE8UNmOCWd29EptB6cP9oy0oGIkd6ulSnHDNonbhizhGJFtFfMrO3NHeR3MbMbZLsb8LNb3T
zzNaruVEIwC3cqBmCqHNGiRr3T9rx5WjAPYhJVjq6UY1bWqv08XA4VMIn0D84Si4sFXyut60QMPz
ANrXGMMXKv1LXWYYb8aruivKXuEM9ptx/vQg3KCEzZ8fTznK0dCfYtEL29+2kwovFqLfhtsUwgNt
h2/z74dXcd7bKn9g2cRNxGpkvabCV8ZW2F8sfiG1Sic5egLw3atJmVtYkESlfx2Sa3JhruI86ylH
MaSPAaFy6s2CMg/EZLkAq7mxt8KqfG40SPDhxDv2ii5q2l4xzaGGKiAGy1lg45d7kuhlc51hxR63
6+7PL157UNChiMgQpMBJFiB14/H1heiWzhg7tA+Jq8mPyyyT6A1ifc3qa9mT509MtSUx6nfs5rvp
+GIiQ4FGZcD8veGWptRIFHAO8TyePojSvqEBZIjKcnIsIfswdU654tKRp6nE5gnCZO4je+9pheaK
eriGYfi7SJLdC37ZREKQIod/HJsJ8/3aTvKIZIp+wDukQbLLC6t2Z6icMwHHOJdwGY1Gl49oSjVR
eKxQxdPUKn6LQjXWRyPyib8bZ1U6d/GZV1GDzXXWKZgm1etAXjLHy3JcGHV9TH3COGJ9AJbGSHSd
vK7WJu3pYIxbwN4o4VDC+rzM6gesnenqXcqWtpqcNclk+/lWrIIh+/WlKhHfvGWHs2vO4wEVmszQ
GKAZCFIx0f+MGsM6aKBFrxQjTKDsWdIgNeNXv/McLs2ro9EE0qm9PysrQqvDlMhGLjz1Y0wkxA98
7VvUHHBdbvgp1ELnd2Ss20iEWLZvouibxlCU8wiamLIUk0vScax4zGc9z+Qv3rnVr7rdAhgYmkM1
nLW0g2RzbvDlz4U9LEm4rCT2eLsf17IShbwla9ZOJsV//owy5pVnjt5waw+dHxhS1X7XX9M3WJBt
XpnuPm389ujZrGqmUSsRzv3GVmblHJ4g4cXgODzfiWe3lu0p2Gx+DMK62n4UMrmXf7+aM3JlziNl
s8BXwL46+vJn5pjXwg08BSUF0sRtGDDFUYvErLGWUnIwZpUeAkPXirFEcXjvj2qZxe3FzRBmhetu
GAQnEujOSiVb3OLw4St+K/B51h3mAzEa57nOPiePYil3raUU+q9O4Z0mYn0Sz/b1pE8gzbsmbEna
Qo8N2o7/XKObf3goF+VvWC+Kmf/lJpwTx5675RlDwfnh91ipSWZiOJnn0KXIb+eCUr5GIKrlE2gG
7u0Z3MXQqXm0FkaKGR9Gf5gXq3locJrwyqE5/OJ8yTIVi75z/mLZdzyMPqKKJs7+8pfcVOTDaqqR
4Zeq0NWEXYn8i0y/mcoOPmwZNw7qAZNhOEPxd1Znnnj8OOwSVoieuri8sUIhYQoL0Ukd0mS23g61
vK6g96oFjgPqkJJpPEAJ5Ajkahz0RCmyTdwGAT8Bbl1cvBsGkL5BY2ziVz5PaqQWf4KVGK31kfop
No0VJb7of3vuISmknJkQRsBlysCwShbvkPtw35mEjCqgObHBz1a/OoIJQNUegMLlYcyef2Ft0XU9
sAmvMuOCKpC53ySzR8sQWfayu6sdNsoDK5hDePKUqeTmOs8wV+BfJOHSLS3mVcZoJ0Up/3glReGq
V88YGEIgW+mbbeZWI8LES+XLlOoRib3uh+CftPQQhb48Ct9ym134AJLSsq4LYsQJ1QKJU2xNe8fO
mDvHTLx+Mx5qWVaxeUo2RLHsL5JxEN97D7eEdiOeARreYgc4JCFOFRskIZ5GvNICYpSA3lU5Y1xc
vJNtaOQXzSGLe3rZj/0ZzBwf+LEjKPtToiaVbwZ2jqMLk01y6UP9yVIuFsR42qxQLX9CuJ0oinyI
e5qZM8vTKisGvUmPSRjDITRcLGiQQ3dDQLgh8PTv7696KkudMeCPgX3QSMqYY5nG/xjDBXE/EC6E
wl5qwCyKX5VTEyxiWRql6SOU/c78OXC9BmZUbCHpM690WX689EnLFKLwxCREFvFZXFPVNgHlJX5Z
dZ0K1P5GClPB1RYRZvp8cdS9zbZPWX/yRaRGUbT8Us95tjmgvy+swWvpNYDPspEWlh82JD9C6gHG
bWR2mGhI5hsFJ2/T+OU/UYbPNbnNZrExRQsXpRXYDcCwgi+Rrh/9F6a8RpNzlR1yCS2SxjdxgKHq
eNcE02nOJkVbGotxscD/uwnjYFO9pSfNZ5cVt4A6kmT+rS9tQdlkPsE+HXoHVWn1MTcNN3ONtaLW
8M7ZUB+Zjy3/riG1us+LuJwtrfuo7g0ZqO7OZsY9KEW2Rnr1jjjyqqhdw1326gaI69pyqKZ8giMT
VzQWPncmCOqPPPEjz7j+MSotCOyGCnjVrzF0ZIdJRiJMrwFIxROcl3Su2taD9vwetmymRnJMHCv4
nXB/apfQ2XPbRfm1koTJrFYQpu7JuZ5Ctx13dyv3JkGImDZKPeRUunCLQw62nA66TCvW0axwoAgF
BF/+H7fqg2oZ9I7wsmWX6aTnnbJLbLGxiNX7oAOKItwBPrisjH1BjbdwQxpnHXUV6lvHbZkfD8Cj
G/5wFstYtylM6Q6g/ggYmenK4tIq4XPlAwq/YSUl3Rn9zIsUedKWJ715QR/YMuLB6BkS8fkT2h9L
PVL+P8hGVpMLfMSnQl9KtJvinPIXMYUEHc12b/iB8MSAHxvllqBK4E197VkZqEB4owHzr1ec8hmI
AJ0Nvvv+iQbg31YACx6rga3UpLudZEuaIkm+UfgV3RUrWo52XEwybp5yNyP5qrbO4fqIFQX+KqEp
HuRe1fk7d/XcC8j/PfAobtrIktHHMOb6pXtJZSwc0XoCWLbPscSCYxWgNMtj4Sr8KdUpl94tTKkR
E2oPPb0K/Z4ho1MqDB6+GoZ8kKdwTbpVJCxruXcPx8cArGw9o+fFn3Djrd9O5icAdLkP7qFt9iIs
6P/bJkocHYhs4bGDPMFmwyYWV5Mz3jAMIWFqxGxl/NlLO/KNx8ZhZke1l9LLGvs24YDHK5mr60wD
dxke6LfgLTk3AfJ9Wsqe+e1CpUdh5SCTkhYb+kbWqTgUCssPjzMy/IGgDxMGygZJT7xw+1VExPyX
AeNsd27YA6MH6J2f8lAOAJHFrg9FK/i1WkbLCJZq1rltNzTdYcKXrHtbuysTAVbJp2TisP2aDzgA
SsZvTVSrzEFUE3OMhKJNGjoMsjiwpQZ23yWVBYaBa/4M2xfOS0D3LVmwIDYtdEc/HDpXeLRBLkJb
fZkyt3myQrH2P6qwRSWN6vyIqzRYXTrhCadGp822BggvrZB9RoqRc2UmQ/bo1v2c4us+NM/NDmEM
GoVhjG7rPrB7vKGvzXn9OH3257/LWyj0eHKGKKlkx9SxsOAuwsZCYPsWXFCk2x4I34t6PNJfwLrp
tIScQEN/HA2+F7hYYCog8XiQheYvd/9yRs5SqTNdM5Hz3YrJCp6e929Sl0Ee8/npHTiOJnyA6GbM
pPrZbEYUye1kiAct0f+7RiuQi5FQz8pbLKiZb2/+EVHakNUfixFrY+TNH/GYdKNdG7UmQxtAX7p5
U98cKXSTRzKRFwEVJRrn47MairojkISF0hMCWEbwvrquDGEl5JxYNFOWxVD5dwx7iEX/e7zRLyok
SmFJfuJG6tUyz2vCbUIPMwq6FUldBbgiYMGTrM/WAdoCsU4RNLNFOxnuX8ijhc1LuTSVrl/uKB4I
ad+dV1yphuMHNoLaoJzdsgOGjZrQg0HJR/cM3DdqThh8pEbv8Qr9TsqNc6ppGMx+2UYXCTcojGz7
Iz4p+qc67ct9mctv3FafAzIIMN/z1Fn4ncSeJ2SqNIlsCAEW7Y6yXTlA8ViXLoPk+NMHePgga927
Wqe24NUzAkSUkAC/i7+XA+RSaq8hohDwUoldZJbt526v4upbIPgVTmJJulIg4qhrC4QCIBoC0UpJ
EfHkzwYua+BrnkBMvGYImG+nMuhvnIXhsokpgB+KMXPdysbpIPn7db7hGFVqZhTlgp+ORFBtTuml
sTcduf/ddF+pNUw7ObwdFXST7FR4fp7O5ZV9tlOeqBQQ6hxnAYH8gOcaeJiCdmq/iGiMhf/GHemO
t2HlRt2ypv7rsBq/PanbFyovULwiIiQ5KxX4ODUd6Va26Te7TFIn1wFVXJ+q158hWGKvqyF7c2tu
SQZE1DI3v1oA3bWMDVN91R83F9O8c878U/hxGRHgYELKonhf+c0I4wJmg8iYV2Ljpq0PBDpF18rb
IwlQ6elYBgYL/pceO92vpn2EA1LUV0Pq8LCNXAotIpvDy/5YRoDR15phlkO4qGJDmBmj2o5gxk7h
8cHdKtq9agDzFZl4qWtMlaeZtyk/kLAT62wE6rEo3iZR9aSmPGYFQYlM8CvYwIUIm+GcoO+pb4WZ
yWCZ/eAnXA0nm9OX2RBihPuUCSpTXxdCJvv3clKSOHRqKZqw1TzhBedDx8s+tO2Gk2eOKnVToTwA
ZNB6CksUVWEhi8HilbckEkpEUp9D3kTB7/zvubzcTyazm9L3w5XgGf2jz7xsUQiWmi8wRhaSy3lK
XRan8YxwPCocj006Arh4T+MuJgMQ8MfbYQZfUU4BsmcbWnIpADq2WfL0LG3XLrDe5RTfNwH49wQ5
r+fgrXQ1b/P+Pkk3ZskpHAp2GfLEgXaInJw766YGGQQ3396O8j+P4OMMSl7m6z8UpPlWug5FZXHw
NG5AVVoWpif0EErmnhogmnCP8VEYDRKlN9NlbXnrKpF6gW84BaeAUgBlwj1jLqpo3wec5yH0KzDl
m5sCPmjadxDTeXfxeeiOIAUjjiz2B+9GoBRfcKjfelN+T+mSTyQWyOsmKNnhZ5DVmQ3zYSLmgSz5
BIguZO2DjCCFFd3Dnxp9oTD/DBKRt68u6+cCxHD0t5dLC2ZXv2eKgCq+1B8HYhZ4ZOct4onOx0z1
1uuJy2cy7wfyroxImU5ZCvcPXzJqhh5Rdipgv4DXD/+49w5+Z2XQruHVVhiizMLOeBKlJRDBBvL0
sPpdj8X9MS4QIlNhbLTBwqo1eCfSkdrXsiWw5aD1pxi4ArvTItzVGW7SAvO71M5XlhLsiBPXSCtF
ldiEOsd69yYXGVkCfSzeR7aszF80b9Wa7RKG2uVT16f206G1AmqMLOkRuJ+Pz4/0uvgsas3rYw28
Gi9+wTzsK9wyBZyjMM6aAKnyGtANnRmzK2FFK2kgNgDmTxVhiNhDuuk3DjiVkNHl4hAFkmd9loQh
ajeUrlbnuWDAGbw8+fOtVbcoGj07HrUHzklntalPCtP4ebVzHZ0v4XkMvPEB9kBY+1UMDLRyLKzN
Oq7BMYT5bPYJPt68EO0vICqRxCasRdL+FSzKp6snH82FSgGFS8iDVixzHRYSLM68V2UXx6yhXCXk
AUTKaETJ4hKhjb4gqBE4rsWK6gg94NNMViKPT6YGDVLKh9pIT5KT4OREMrWoJmprm8rNOZp2sfDT
D/vpVT2+vrxXql6kWXXF4SC46DtAeA9m3x5lglbRCY8RVO20R0RqerJmpEdeQRt3grMJ2YCXlDU3
Fax6l2rPT3pRl17gppyVTim5DwDHivvwQBFxxdM1i+smMAwOwGu+pCX6+chPsrvTH/UReyFJrOE3
1lXszUuRL+3k4sqmfNM5n43+mwBPI3XGwaMEkrqiKmm1PRivgjCm5gibUjXFqZtk6d0qdFcyHkoa
Nj0L7we6+q/oFMuZsKIFMX1RL4nAgmf0RQ+Ig88R6hdjYm/KRdA3CAxsHQUSYcZg5kMKxuIe/D8/
Yfh4V1dcsp7vVy6Xh9yrhjfPVbqm4AjhBQGwHre1V11Ja0PpW0Opi0ZrFEf2q8F/HR3w899Tlygl
iW9bFsUCrt1DCRgoOeS40Rjah+DSKJdNjcjYO7UbJYGkM9XlHl2Lh+Kqz9/5IQNMUK+VbQFdsi22
Mkq0xbemR+uGXiqx9pftxejJrCGSJ0LF3Xt2ot6ImmN/Nk0Fwsp/0BlHvErO6WOfI8GSCsN/hEsO
oelKTRxIqWwv8ehGSXxDuJBg3KS1yfq9uTkcOn4QlRdtQ3VpLluw9/UEdDDw4LIP41tqutog5Hy4
uVPrptiG+O9fLk+5p2hoUlGDHHuFUjk1aMYCne6+UrQbgkWVEcc0AnMpn/GcpelPp4jWZ5b4kH+n
tOVpfWCUbxjuJ+iW92d/GtIpAUC0m4cDW0PZWc7kxDxe5On1Aej65swHa6NVFf9eBRy8KRjUlL3h
RehUwRbrTvhnmQwSQd19yG8yb/aKvOe3rkEC8U6oVe1W4htL46Gwt8a1J6XYxcZf1Yj11CHGl6S6
IZ2AKJIrW92J4gchSASPuK2SzOyp1ghvHrXtMb5pQvlYjevqK1OXKu8UXDUuBscsPWZgP4AeW/R4
0f2FBAPoJMxgZ5hVTgkV/5ItnLttgYB45g6AcAc6ofMKl0t8mxxsq3m3IS3dZHhTre9pfXbCnuWk
nafWSneRB6WR5QQRRH3CHpgEhk2nQCe04fekBN4EgyExIE5sy0/2/gOdXPQTYL1NPJZgCo4KUgPQ
N52DGn/9ttzUCSeJxZEemGHv0o1MewaY1T+9eRA7CZuu0BYtBzHgOIquXcPsA9TFI/JfYFP1uaCj
8PjXN5y+xVJnO42LRAlWAnOLSAn31JOwvDomWG4N0Uel37JoHL+dnuNq3jmGQknaoAq4IFZYPcfq
KgZtAorXOIs6hnOA3OgFWAq5ddvvlUcQhIOE/jg7drszTJ77DUMuNR4u/lRzs/k6kNAWeXHhV5KS
f2bUrHxXNnFnJx7U62464VthGfYtGqmf6DVyO3zgfs7Nx/RoU+nv4JiQiRnQoPG7XHz2cXlsUDmc
fQRE4ukJycohwL0ieskNZ9fkpEE3tbPGu6xCaQ7Bvh1Csx293BOi/UW0PelDRW2fFw6Dy3v8s/7u
4F7e/1z7wQPr33cG0+YSgl7m2Eu0zKzT8NjSz1zsmHNaP81uvCXgZWCmsX9YoO8TVfP9r1iMp4Xx
fK25YX+f2zsHdCHF+rzuj+Cr8zXObB5OT0obi/jmaY1QrQHKMYTMShCZyHt8cDEyDqPxB7DZ6Qd6
8SSfxHvWr22MpRBagdJxSy1Z+NXded1q6bWS9Boiu+TxyX53dUVS/3nEjeWvPqSUGLCq866xndQ7
qrdOpVqxoT93jFIRlvlnH77dEPfLcD0DfYIQsmRyFgzhedDbLTMlT5W+K1/tLqYUQn6nYDOSl57J
V14WoICch/2EOHfBeOzLDepnF/u01tDORahgCyO73/DWgr3sgwqLr6ZA0CCNUoXGQmR9wUI6xr9c
Ig48MfqBd2CHyFzmojKuiLj4EQ2LbkAT6Ucnxl/L7bu7shkQDARZo4mvuedekDH9xngKXSIsbiS+
e/z4UEKGKt6ph3+1/2/w2EeYphOHz0sXZhSL4amjwc2BChVQkHd2dKK+jkmllMRv4HFfmRfXXTrS
mYu0SQdI1jkTTqp9muwgZXFObXx/FWKOTQG/AKOqDX6X4LsMqWUHak/ucr39+bDJZtiFOtgEtgAS
FZUxAzYtfM6L4j+N7GCDU+RqyFtWVKmbaWHTrlrqhWZNzAT4vF/7VnjkVaqWjhQ6WgbcUIK/w09I
F32bMusqxv4qUbLHLhChM7sW4d5140etyV+w6JiDhz8LoDe8TelznMEmv8LZU0Un/ER38ptx7TSM
KzqIULvEUAstvuUkSUi/e/8mrh+DQScju7fPbgb4rrl/w/BomLvt7yqzWdyrFkREzpqhuwNpGx9V
5J94Ex0dFJnBo9+1rQQ06dBKqjmQcy1q41lVH57xDUppeDniynM2JeuODe1m6TRz2PwdeZGRjs+J
kXn5WPEqOkYL8du+/30kjcSF4RPUYkLKjoakbFH+s+JXI8XuCMIr5ST27eKBjxCQZpX2wvB1TGdS
LhHjbDaJl1iKWMP7RegKNSqe7PS9sKlkovCk6oIOamm+wcbq0KHkXr7Lc34diKzxer1uGATPaTyp
+fR/dnOVvoDxnHAU7wrBB52VtsD5YlgFlK8/n9JWuGjiUdPnZvG35+uuCaK+rdtuD/3QWqvjKe5n
pE2Y/TU6pKPjpL/QqInBmIZ3DdJFIAyyEt7JgGWItk0OSRSHUzDqgEDDPhpOxZ1tV1cIqHlGVWBe
1zCcUp3JA/oiix9FWhIpN0RNO88aD404YtvlxaB8SZSc5o3k3OgGld6XXrhxtLxBIlh941cP/trN
TRXFi85hWdr2Ms1G8LxsuXvI/mK3JRqUoscZc3RQeLpUtnZobEtZC7QJ11iMbyiI9SJ9y8i+6qs7
Agxt4k+7Q1UWlD8q34OMM8GBLKPGgT2ucaztzklSrTqWtm3QpSKmQS4Z0sg2raIMdV4uQTkjPhR0
4F7zxkxO+BBnXggxSnxZbQSJosHpOiCkat2m5jF/Pr9QWMLGzBrDEOgCodO09jNwY3cI8n8lSq7S
UbNQdmlWrQ95o4A0liHw2CT6apoTSG5eAzBx9oKlji8T0RdbnDlKCL7VcVjyuoD18ZTKiAP105ud
WGx76nPY4wGuauRJydX7i+I+fJo+9CxhhS6fZyJncZH3RbUVgkyVfm1Fsu4en0pTB0lX/nPPf7i8
JyG41DtHw75BkgnYi2O79gJC7sKXeZdK200aD/3y70a/jg468XKQGddHJMD66CrB5aenKGOr5KYv
PUmoqelkbS3G3d5Ql4CHDniP0my2h5yLHbRSFkRzoz43pp7y74x8fHJqyaO5TOLCKSnTmPh0wk0K
kIOfrjo5B30RQFmCu9n0uJf96qcYZWQX58vj1I08CVE4IPsl9coaU9wf+HuZrbTszQi8Lng946LQ
IwB5rNPETJAG83LgUJbvz8fZX6ijFwG9fd8oj6w5JX4V+P7wABNLn6AlT1MG4VEK6BJlSZjGTc0i
q5C3zXsvNqMNSMpU93ZByZcjKDwhoUGEmzN6kRpbjFaOvhdsuMq/AEPFhR4qpRxnpH5aore1Q69J
08ZnPZJneqHSItomN0bmfGOHyVLyFBR2rWZPc53NQF6mnSTUzFCd9Pxy+Gy2rfC6b9uHFT4CxYNt
2zQW8bqP0qUGwpeUvZMSj4zd9NhzNVWerlFNqYZ3cXH/x9QT4+TxBLylwxWv3vA400gtcfUOtd6V
ylRkzhr1ymCfV4gAEGIbilatWNoHrpRExK7bX2ne+g8sNTX+2+fO9PCAwLq1Y0WZ1sivVPFvILw4
PbDZGSiy9F6+NOijYrXF0m78uGVLOBo/i+ZPRxaJHd+ZPuUyqDqetXUom6i6/o13rSe8d3Qb+u+C
/d6DRfOgVHfysHfh0Y3AjmEI3FlrFR7Y27odv/xDB51qFYKAzw5H+yCLv6i75duh8NEsFxGWfL+c
OAkuI3eVjwPmOhCc2cJxYxcekPWNXbnL2CulkAspr43Nv3HrGhTI31aL8J4GND+VSgekoeSpo+wB
ZhEali/Fs5TupQGpF6/bjJeRK8OLpu16rqL8lJKIqWnFZq+5YEq2AIDgS7TN2TiQDIZeeqjE9PpW
0aueEUnTF9ZUGLUNYWiTv5AJLOPg91wl0C1GnhwB9tczpTruhzOopX3jKug8DbZefRDS4BQJctn4
PSxRdkVWMwr/IJQeoPZXfYRcxWToIrs/vq640DnFhGkOogATRlTZaTKG/dX5mrInNHNFBlf2NDvj
4OYt8Jvj+p3Jev6m0SGuuRlOcauHbEFKPbkPMJcPv0EXKRMjHwgVUZZe2Y04ZIit05mYa30s2rWg
+Q4KWejwAimDTwGCKStu0hB4rs8PeLwu90rPvUigd8+3uKHxy1n/RSFC7rhRrmRmC8Yk8kUenT5K
9E6DRnI4Y+Crr3e55dNVqrvDzf0fhmYkzbqD6s/8UOcHi8V6yZBIPhBpZLdZpNnOXlHYI04fhZqL
1u3ktflHoAdGyTGrWG7JLx7O0RmauHooypz7NJNQU4plXg1TBfupLN1Qsx/BHsrIDD7ryY+Pb+fk
pIt6PMN/mFN+TTC8WP9mtq29LmU5o3y3+Ra29lGzhjOlAwigp/R7Xrk1V+pW7sHhPZVGHm9Ls2r0
UiXT2aFVBAFf2oOXtheaMjozimJ/+428IJm1D1HOopYwXbVbEUetvOPfXmTwnrvWE1lne72wLjxr
8C4A3QBbFy8BWsqLR72b39oryh9d9B1S6TRnOrZ9c2MCcJeGGqZc9lrzXSwFsYeEZZ2dYRFnjGNy
iyNlnrieXcmVjBCrFxvAC6KvX1uWZE/wwsPO1JW3GVutZouEBnTy45HxIuoXhCgdWyISUqV2krH1
15bnDf5LoIBPVBPyXnnR6Y/F2Y9qvsPwrLI9fF9V3oMXMCpXBeeDh5EP0ooUNV+ER6V37T/8gPyx
wDwo1hxbGI2Dg7F+RB66jsPbWkRstdkE0k61WBM4frnTdv5twvmkWvBqI2IrsQWPMJmSUN+/wX3g
4EXx3IncymUvcacVlUpmplgQvZ24TVJeAlkrWFZyBj0HVxdqHxh5aTt2mDfFWkB8rOSN7NI15Bdw
uBSmZU9mCBPatlTUx8ba9+BbUuKyd1sd98pwhJU8EWyygEXvC4T8AldiA0GAcpXzy0UIBEOfjbgI
cwA+A49FBuT50bbtCwx3Q1D1KAFuS9vDhi8djLQCWFNQAbKgdWf66Nh6Y1DFzzhm1R5/mxulb86T
5Hxh7taym+uwpqssfHcJ4UMdy7hO8zrjVhYLcRskxTdbwb+55ep7ns0ozfaVkZ/23geB2HDY0EaR
Imawipqfck7Q7hF1/xjXi5pGaPf76aFBAOyIL46qtINf8NR00lQ4jC1C02V+N2OR5QpyydWXCXJK
BC3A737RNwLeG75w3lTagFtPM09Cv36h4ZLSwLxVkvSWlCb4BGVqXROyL88GmM7s2rMbsKLE8SS6
rZAQ/4l3bsRxfkzKm8TKBSqZ6kLiIZ5m79Q5dJddMgsdYImYrQsFYHDzLmfElS8ffJi4Y/YFNhZc
nhixhEd4F+OCyFEyXzieK3DURhdxSr7xGrX3Ymfv5tYJ/FvUCwDqNlhoLrrjPK6EsJWZsB+S3vvz
Sp7SOBh4S/e71mT4mNCLUIHpesnTadeNJRFsbMOz11Qpn1502V6SpAflN2WB9xJUHVtDr0oy34tc
XqAy9BEcEG7/2fOlM+XT+8to6ZaJZpyqqL7saD5ehggQo+Gk8XbOvFp6eTINnKcYFIR2MRyOC9/e
HbIHUqOHIE9/13BZ3cTEKAuA9zgRzYcSdyH9/lm4xXF82E/Ff7Dol2bwnfaB8W919ainYIVvT1iI
qs4bkUWTSfIDMGd72NotADanAT2ExRAT92jSgJpKR40HYX+RoncDw7wdyh6Egg6CqRlbVkL4H1zQ
0PURtzK0KpmYF1vdjMBN56oPybwf83eOhP0DB2WyE4pw0oDcUKtpL0JqE4rYuZwLolKZDJ1IqzvR
Ap2RHikLhb9t+jK/ogCHjAm5aeAOEboG5IV+h4Jwy0QAgloK3nkTWqm8SBXE3jKpVe2HAykieAKT
bgJEM/4ukbxLoInK15gIAyefopSoYfCXsNcFdZSFnlaiG7cu/kd0gPHZqUw8utVkAw5T8o0+d2iP
yYs/ArqzmciwQ+dyFQoXS4NZ1CHI7fzoiO5GSqP3dVKP1acFH2rPXiM6nr/u+QbAGTa2PhWSp4DS
9gp38TDLyvg0rJmKCvJHovOJJV8pep96oDRq+3kML+5OL3HbCeSVhKpnsHbTHP1IrEUyhOy56XHZ
2ztA1XkK6wzpmHV7L0LySnNDOu2FuCNlWA8PHQ3i12szRufQiFnzrGlmAXX2pgBb/FpnUWd1DGDb
avN9c0T+yCqfHMl1kaNA0CQKr1j65VurHPFneipkgDhLxz2upsUdl0nbbBz7f6s7+YRBlCNQ2pBj
7X1PB3Q17bJR0hSiHJiviu6ge2eD4Fp1g3fzs8A47LIIPyPMP4q48HAMiJSNDAEVP/872G1/tdyr
Ib52TauLlvbf7+3ZvRJ1fWoQ8YfuQR5X15iTSyf8VXYRM9BBOk4eLtgmBbkIDN+WlaMBQxVvDfk+
mNLsSplnL/uGTDdXq+Uc15cUXnGDTgCkiTbn04tPsISkCenU9CcjATBeDj3hBfIIJBwcCm0gbOIv
fIrqUTPuG8TRkeZZ8OXxw8qaNmNgM2AeniFUGcbBkYQIxpYVeVkkX2NAofErcVMiGaWqMeS+7nhm
XT6Paw2M+Hmmj2EnRu+uXx4SPcGcueP3hAvU4VX7MMfeOTZKcVJEWOlbCA8hrR5WUwMKyz3cH8BC
D6YnMPoKiBgNVS3Yhegps5QXoDb1zdjeA8QcswrOraPhsUoE8P/APxdYahtlnCHluhAYquhgGUcX
JAIhHMxYnmJQ3OvPhYOAU+wce2qGdFFOdFu1vI5SSFKkae044Vor1yZUCXpJAUiwt7Fk+eotIFS8
6luCNfDn3UN26coZqzqosQ4mK5n0sjTTcRUFgJ/RlU5B9zxYgt0BFvc0pKEIcCNhkRLou3e+tFLh
DfhmZP4zNX3jlZIJIMcy1GtldSzC62n6DVMwag3qT7nshSP80o6oakMtQ6EkCuO+sRx3Sg6nB601
EJA52xw04ci5nM6x/NTQX2FqwzUjRLrrILhJcFKg/5Feh9owhzRLBacyVyjy750/Es+0zNUiec4X
1VzxlnFOqNG9hDbCHpWKz4WwMfNlyntItt9wGHrHKBfmikmLl7RhQTXtjcsY/yVe/GOPgsYNmkgI
mkHAkDoj8NPD77Ni55Dcl66nxbXVs5ZJU3lumJGVvR4U4SZtoi66OdfB0IODHiyjxP2g6zjvbo3n
WKDFABJrPbRbCkAY9Jn5dFe84msCnYqgH6l8nnhvBnH68ZKX0BmfL9dOeKS1Y5XL4C/iYpmFLePR
lY/F8xfvcpcKspoohH1jqOKdKb8TXyfb2b9CekOaSscQ6u2azdpNpanJjI8Fn8jl9fI2lrrCXCMx
IgGhvUfVFay6iX52ftMq05/rEVCdjg5jA9jJLGzw7GokatTIrW6w4sjLdvJuoNPiZDEK2nYjZyci
pSimmwE9AEghWw435s4DOFgRlxJ5oEOVk6Zx2IsMvk4nk0jz1sUSiK2wqQo5W3OM5qLrI6rtF6hJ
GQT7nnYXQ+xKkFTzxmJ4Cx7jogjpX9dq2wXi1TO87A6eWy2wUpX3mi2ni7yOhTKWVL4Jg6ehNE34
9IZeHUgF5Q+J1+xVLeYAvxF9sYWcBL2Q6GOE5IUZ1n3Y9iuaZJOe3Ok0AGnQJppbOU3ed0JSHJw0
M/VqYwrU9QpkHBY/6TwC06SyTeCjTfQjxpIvVISlIgGw9U+67fmh6Rs/8PfyWKiJJgKNad0IDkDx
XwiJhmdWvkIjHZW/HvQiIiPrzgvz3sschRRz0xIbgs/VRfIUcfI/Zzcq9rvFSB1sGmOGFZTMLCgL
Q6xkKbhgRMVJH93KJltFHo8nVqLr0X695iHm0aMZeiIytrzmqYNtu4KTR0TkyJ4VFSSvxBGrjPw/
V1g7IW/JAo1HYTRBhajwmNfB20GXm1xVH5G6FCSvctKmAD4Tjvoq2SmLteRG+lev8aEICLkrm8pg
rHJ4KXz1iIN69xzoMXVIGg2YREkOSA4zpcv7xEAxkq130hzr77cDd+YDGxdWFD7kL/Pps2wiSzRN
QgLGs98lFU4tCeLuuJa/rDoJkSEDyHuoXbjXDhysmWlnNJiXYgbQjJNTfNpFjP5grSOLSQgC5FV4
y1ma1xeqOdveNFEAr2ys9JiUdKDeL/haHGBmViMFskdlOy4QNo7YvAPtS5cHFYjND2VKKxwuaxYR
UGprFkHutKJowkbRS8RDE9Fg729l3RxtXhXlv4JIobUyBGQNnuUq72D3IVz/QyXFGOGFfLvpwarg
X1AH6uqRWJkMZVdHQyvzGgM8qHuSgG/Dr0F21bychcywzsOaozXAdtWU6HuvXCdZlfdWFtt43g1R
h6SrJStP6hNIdloag7vxyrgaMvLMf423dbvSll/mmluaozAlzdYid46qCU1JjIAUM0LL7lYlQrfp
Rt1ZBVYnFUEjyAC0KKBd7wmyNiUgVnHU/Wh1QgCzgfhyQDFCNOpCYWs+/UTwGtF1QQGGHw9UVc8o
vGgYOkNkRN5BroF7QkjsxyWOtLC6MkuwU0vS6MW71EW7CKQkCq2LjCerUowBVhyHfj2qP0MECk0E
U3YI7BKBZbnBj7cSN0HxXvRhCO/v3F7owgRslTMG0A3HDjHKPUyXMpXhCGCT7Bb8vtaPOqfn/VN3
rrxTajJ/Gu9sf6dPMqCBOCERHJMqh265md1hbq9sa628Vl/nJ6HAvmSt7tkY0wfS0aNtGM58QN8j
KmPPhsRJI6adJj7Y51pfxOY1FJIYl2+n2NZgQG5MoibnO0MUBQP39sgX7tjkS1YB/klkvS+BOxYM
YpocT/n4uxpdtvB/XLZqa0Wb1neUqCGkgwhJjXk0KUXfIUUEk6F/25mp7vMOBc9pgaxtR02/HvIv
FDh11EZ6e8DWtO9x6bqppktm5ptctFq6MiuK6nlSRUxACPu7KvgHOUXROgaEjFAgnYQdr8+XMdIO
2kMboiCqMbAFPxczlyQ1Y3/dq7vuFM0aaZSYPDvbvTFxtobTMpNvUzb3oqD8+g6cVgfl0XS1O7CD
h1XGzZTRO5MQPFDT8DeQKKbQWj1wU1msRWjmrEjGcqpzYA+DMwKzXCXI26u5yOQrpfR4wiud8k3v
0DyMvpuPgLPyyRUwezZrq+ejKM1qceqGiqH8fjv5QnrDVE7rQKEy1/RgNPbYrdyNSbq4Ixm08paD
+LUtbGs1t9IbeckSKWAMMOEH9IBqRNaNztJRs5bQ2P3xDiaOkwqNbV3e2ypOFvZNgJVq5CIl67Sn
6axEai6LasQUQd5ZWJNyxrxJataqkMZ1apcOVQm3AQ9WSBmYrO4DXTkvixfU44WIxEh+zxQmuS+t
iy6UfNUhAaBD7+SXwdKwKH1SPBV631icEcK8w31mPVtpA277ZblByLzkJXPBRP2meDovHEves7SU
4XqeErdXXyZsIAvbOg9slSJKe52ADs5FbzV/Saky7TwnFYl/RW8vSA8ejI9xwyFEps+9F5oqQk11
v0oEtB4arpKrEiXCghcR87k+bsoevlFfTnSk+pYZbIqbN2l4AD369t0xFA9F31zVaMveTTkK8YKZ
GKCNPyrhei2VZ3u2V5oSEmWd1QY+30mngGl9jB/hghRvqtKS0KFswgg4kttsxId0ULdDggx3oO/A
6+J4gD2xYt5GHI8tX5SoXr1yKjId7r1ahg543XrW8v9dB9rugZ0nQOmOTCvOn+7PD+HvGhMOdjL4
g3zwlGdb4zxExHu2JhBhRKTaCBH9cy2LrfwHvdke9a4O67zqlWHzGBwB5oU8qfquL74MdM8Uz65G
QMRO0A+azBOaN3wz7nOlItov4HwikRM8cudFl7RXtPZArcJnt/vJks/vvJks3nQ+QB8ChkLHOBXI
HmOxhtAp6F4rAdIvHqj1irwVQZNhuc12prx0qUxR8jorByB+XpukiLelW/5RRulmTX7E9CrNe+ID
4notKOjPR4X9OBLNChfyIu0nMifSMqZ2sElkxVSN3e878ftcnHUhpwLLhc3kImhOzPVXEXMgDPko
wHCte69/WwAxz4FmaKgCkYaqzM7ye5Hr+PC2csw6MePu9bIryctdldl4WUB5hQpLlrvvmPVvJO9g
gDN/Kxkx66h6UQmyCaS5NlOLLEAYsun2yLmjXiR6HTBKQ8QMwqGP/tyyZ7i4Ch30kFPRK+uaSVmz
yGNdGXYFFt7H+s2wPkRMENRqywwFIt1HtlqVclzP+RsZJ9rSGFPGHCaIEwH1eDjLiTXNEGQOrS3h
DdtcoUd/niM2b5GPj/Bq4sP8/o0QMqrvqGcz8fBf6K8k1UTizql0SO2IB/CGwDsv/PJC2SwxkeJi
+/RfisD3LPGFhDxSTJ66a9CsJl2IhZ69W9U/M8DLHGHt0GfCLYu9ZLHrICtUZl9JOg5yutg3V35o
8ikTWakOL+MvDRbdzFvd1nwXUVS9EnqckwO4cGWdb23wChoLfC1pg5Wa5lJprMzICw84lBPveu49
bgAsPCss2gZl6pwsMtItjvCdhxwWu7c98N7vZQnQoV7b9aD1jIgVgazNfedb/vv7ke89JAJlIx/B
w8zHB5X+1zUUaozJoJvhP9mZIz79e2Ur9w+1TmcNiDSavnNnGnDwmBmKv+UMm/0XsFVXVxed+XAp
QFO2AVCN5sXDezZRBkGRZCIXgN++DT4r79m6TokLMWTH6UytIVk/gZzqiUmpRbuH8y3EK2mYUoZN
3YYU7EZKQy0QgLM7KFf4k/nA4RJ5axU4OBMOKVxWj1nriEkerwsTW1lEkxoGVtQf2sHxqcpwYXoM
1zLKiqHpYgErGyjgCxk3fd5VRJ//hXUzf68q8bJzOGK4UizxXDNtkd1ubsLkXJhYzq3BkBczRnHj
wgEi9cR2mFv9UGxAvn+dmwyvKpGlzG3TmM+qXrkQgUtF42CEg9I6zQRWenWB/HcFxrBQuCu2K1DT
yfoqM4gpWLc7CqmlrCQQYWNNfyqxOG8V1I7RCz+2hZHU62Wt/lhNlfLGmW1xMRsMAQernj4Hpmyk
om7LL3HReVu9H2zYWUY1CLls9ZcdKWM7iFQ+r92A1eK9deoJOrGfUxOob1Nfd3aGGdHjBEr0Rr3I
1lXHYBF7prEi5omTZljsJBbWmORwx++o73jXtVH/AWkLRMfgJp3Vq0QPH4xB9v/jRoz3ijyJZsRj
zA6tN9YmrnU2V6YWbTMIYWPdCucMyXyvYU6hd/E1fCWq/AMpRHEeIXhMI1WHneNlTMQs06EhXwqW
eGk95PCKu0LEYsQtOyZI5ujUp0ThttLNIJuOyw7SzKnO/meMBpvmeN0PbC7dbcxnva+c3Id0uz/9
4u54vz7BiiImpsmV4Nndr6NINE2ovWuoe5K6cD/ZGWQNwSooBCAqz/nzARFiP/4Qi2ENZryVNqMq
WQfcCMubWvcATJAvqUlRO9GWnvmK668WnpZTVH20P4RuFh7CCGA14iC2HZpgWUy0LoTTC0PLiZv4
yrzksaQhpeNyFkmzYTuz6uyh9TxCfWHK8XdXs6r/WVhM4Lozlrvkr7EJaZaxTyXWpnQIF7In4XtL
JMxidrEAX8sl9POURIhoDwmEkStAAb+fnolNiMXxt9K7MlU+0r1ZKMSWMjnNiqXzVOHGXsKr+/Ii
RAKR5LhOs6IFMVzUYzqzSRwp3RqMDF9YHk8qy+xPl/AD0ElBAhHsLGEl17jyly8R0jYkvtqtca3B
ldJ3t+ram1WOQrJB8+C3v/qaJr0QT55ScePBqaNAdniNNb9D547G6Kb4iMaPGg14HXvBsaYzLfKK
H47U7l4ryJ7couvQ7dOOmnkwd+36+M5sIxaWKMM2s18XxypSFoT5I1aSFCA9/ti2RAM9zWayooPy
DL0xPTysMQm7lDsWOJ6XaBKG+p5uxcUpjVPAWCe9fFWsLdKjv6QuvCSBkgCzvjaF6Di26K+olcjA
2Y1O88JKIYYj/eJcWW2IKouw1qNboQf0JbMqA/gp+Vl3msSDezptA7Nf8iskEpgtdXxFYA0QEH+D
REFd1nX4kuDi9GL3JGCDELyPRhY8P47y1ldlukyH1c543ldp7O7RY6FZmns8ZHZXSvdzU91N6XOj
qYIZZM1Jc8rVXOxyTJs+qJP1mxfGt8DLRO/VfylW2LGJvHJgI0qPMXy8ahI/FqWg/BRRAUuEyvx3
ZHAnMvItDi07o5Tgv2mXsYJEB6W//pJ4gKBEho2SBBl10X89uMh6z9uiaAAVeOD7RePsX5jYODOM
JNbyDD2LXtd/cFBihCVJAv6TRtb2bWwdAmwvInONY8qiajZzmozsMmokPk8L3y0Yu9oTaiA0fYVF
rApVjvS9sSidT7/5s9h1o7xC/r4aiFnttiEgaHWVXFwL0eQdABfpIIjA3nivpzOCK5imxYcap5PP
gbZ8EBVK0+ri5+vYmYqw4Ili0RLSBzAvHvgHwkEAYOb3HWZfsKjdGIsbDzBD+ccnNDN9uhTOTHDU
6QpoCRjnW+CKGLH9GaKex97yTNnvvLrshPGXD1egJicm02lVLzzp6jhDdyXG21FRiAwofFYmtfxu
XEnx2OSME1HsAdlbnm8k29e8fOcJfvwJCypG6tXY4dXdfYp0tt167PqPsbPwl8GdOPSLIlNcEU2p
VympFjI+Qe/2Dr5x3CWms7NpidMG/wg3HZ8vcvPsqWVU8mWJgaD1/UG2Ixjxnv76LB8ofFG2Jb+b
ayOqoiBdfYcnIemN19KmBVpDMNN1Jy5QMy0IQEoXNHfeVcI727YQwTfT7XptSDORv/o9LTjJ8EjC
fVbYM6V8b50XG7SF3fWMn2uTeunizl4zvKbLsVaeXmfRN8InyZAgklIxK3yj3jeO/+Q0yZoR4l69
/BUjTtpyn3pqevumE+td9ozAz5cms8VmwydcbfdQ9prxgApz8Q4Z8TSv9k6E83SGEbh6oUzEbeAL
2vwhHalkZBCIPcLF2vlz+yCcGVoVi4GboIwPm5XczpesUfhi+1dr9aCIKPKzfYbBCy2mKVzWxSWs
PM7VNh13sCwCaZ0KrZd4k8RWtZ8cuefJ2maPhOVo9mL1hO4+r6QsVFeG4n9ZN9gIZESZpB9xqjPo
opgASZCftIp64qAT/mB5VnF1/gYahv4jm9mQ5v5TbFRY6Wrq7jGK8URPBTomgiz1jJglHy+sUU60
2S4C1OB6WpyiZpZlq6w9hiiNGBrYV92BbWiMQn9DgcSMGTWNX4j4H20UTOvNF/oblXL1Oa4uDJuO
Q8Ylxe8vxlXe9hFP+80XUwZWS7jXZGagyu4Cu7i4lFveOJB9aLDu47V3Bdwj9ToezcuEgcElezQq
N6svx7SDbXbbrQbV8OpfJFFjeRyKgq4TXsfie+BYkcXVSpzUKjjonvzgS5fp2ak6iZWxsyq0g5Gw
fw0wuceN/CaGcXtWwzM1v6IjAb5/fLiZnBz/hRhB+Jnx30lvJPGfQNl7DCpSWX/iKNppHq9Xjx+Q
01A3YTDIkLZImYvFouRG4gWYQJYMqAx5Nb4iQbHZRBP+AizvSyumr56SmM89MNkkYPsD6wG6j+CL
QWdd0d8k+VDgbW9nEAeu+CwlJsA+DDkBonLbk/zBZkFGtNDQvA3WzDUhlyGG7zQQW9Lsdl9KAVw0
HpeHy1v/6hhsnppnxMoiWtdiW9+xqehBCMKx8tmEFvWj4/0TJIMG7Wm3Wtfl0U/L6epcnA6izAxO
j28RsBqpI1EhTRwrtF695RnR16+bITUVdCmCUt34Cv2bxmxc3K5wA38RlIUYZlRZOjVyeSzh7LZO
F4AfcOlvYrs1bmc1YK4NW/Y6uSPEVeW59A4VKkhyAE6ZfBY81F4vN3oaPBhDhEt5vSLfIybWPFW6
0IQXsrakru+e8nAbcA/jFQHPRMDld3JxYd94eYzjXKueP/wD6WjRKpOaLAfC9iOzrAeq+OKns4m7
nhwRTSIhlPDYj1YU7ji+kaPd5bTJ7/KhL3d7ETi+sUxuEk/GcpxzYXq8GSjb6UsnROd8qWDYH4ZJ
3jwb9hwjLQ2vGRRoWyMmHzvR4bh3BC66qFQiT5K1q3z2JbJtvWTUZ2phBB4g/EqaaDQqrpaZNbOL
3VTLfa9TIZUgA7t/0jtLuJ0NvYFUB/Czg6pn1DyhTiMgKaajsefHM8bIukGQpHd4wL7IdEx2Z6ma
miZhdyhWnqOQTLwZk8E5VLYShjp98dzkwly2+Mjo7mUXj8HyYJO0CP8QM7lBlYWme0zVVIkuftN/
lRuN5GUdRUr2322zSebcNmCfraosa8/EMFb3eL1+d36H06RxgO1XoVsSQ2owuSk0ApJAXdMjD7xH
Ualv+P4env2k003pfFa0EEaNq3d/GOYfgV9oy6Ae8cmeCUfyeyRiKG667zvysrZngouwQs8IlWvM
UP4SqKk+5inyOWtJSkkKEikoiecly3myBrhqa7jcHVcbUr27xlRHxrxEHCiX5tW0tnnwd/uvNBNV
FUG0Qt6SQXSCc+2mjqoTQWOcq1R3GTA2XVQZmZTl4W+pvl+zmG6bEl4sqrW5sa2h8P1+FgI7EMtw
CozwZm3dhxXmm5XqIWEYUjRpmwHS+rsaNecfKlMATqVs4y9OuwmckowwoqSTvFCO8Unmz4J86itc
jGcHrIAwauVLvznSyLyzAEiUk4zkKqGvSP6A2Wbk77yKClalGY4oCttYv4exIZ5SNVCOZpdUC9y9
A8zYi0e928WP9DFdoW02Yi6cOyHqiubTgqT9KXQSwXEzpQx+z8UvPNYoZPHUkAR70EotAwRbzp9l
0d6EsMbRw39sgkp0nN9dgC9nBtViuEZwFqvenMsGAxTYuKJGNUNyGssOmjyCchXfKZUJTVWSKuaL
oFCspCMTC17QdkeujkpxTvRIx/9Z2gqcFjt9UUKZcXy/CUuPiDUIj6tiwrUY9uBFKuQ88bR8U+Pv
FQ5Mbx1/SNdXiaE2kuK7k2fwKSZ+nw8qc73xd+rcMa/eEG7GTVaxa/vDnoldiuDP5dxndaWew6lQ
SjkeXmiQkMQAsK/pFJzg9eBqL7yTOz5bMrbW3kjqL6q/toVP3RO4CcJphn1LZ0i7XhfY1b0sobsE
ApZgJoGEl1tfz/EW0ZbeG5HRpSUNuw0rm2NCRUllgZrouzWA9rXcPJVbuCWa57auxHCwGaZwoV+r
G/CCLG24Xy9Q4rTdx6vX1DatuOGdwyijcJLhheZJoU3r3m4s1Niu+eR8nWITAKAEpD5enKETokM3
H1YRZ5t3dz12ONrFf1m4A7PYZeLwp+7G3S211XN9qrdKUXwhl75FxCDtfx1NQWIKmu3GGjcYshT+
+Gmg1jw8i5lYHMewOwq4HsxBOFbGBWK6QrTpXhXr5LOCe0eucahzc6exyysMdulx5why3T4zcATK
xfBnki1wVvQF26afjKMX3hPTWWnyRfBDbZVeiSNt1nlg+l0jrxkx6hNF/0f6doa1vM54VVCbK8jc
Att6wWErAC0Zbkx2MLNRrsHosIRw2dqNWQkALj7ZRkI1PR5+ObmnaXv5cYuCSDw+K+Dm8024cWYq
KFljnGO8khJ1mIdI/n+uy5bmyN+fXa5hb7EuqJ0dKu3jWlpKNAn35EAyxQTCFa3N5adtaysV8H6m
+7kz8rCyb0QOWMg+ji4PpKXhJmbXqfKqE7INBSnOQUP47tioIBYdCNSw8kvNgGplkTQ0/CdZvHJd
B8ENYNbKm+CUI6PkA/Ml3pZcNo8Bq/M+pkfUdsXpaKsg4Bi19ggZCQ/AmvQznfbA6oUEB0WL4bYH
QYWEFK0G4OG3himX3VGxMlpQxurOHKL1qtkRJFFGQ7pjc5F1OZ1AuopAobJInFfJzAo3PuaD7buH
76f8c/6WcrLzgF/xlsOQGbFoRacPtyqqiTdsLhQluUx7ktbzWZ3hGxE6qQuHFXOWGBuYaRC2fnkh
Iepu1cloFmAJgda5A40sbWblyWLQx/BE1Ec5RgmpLsi1gOg2tDAfaiY/lq6Xt3ROVM7NbeVONVPJ
V21uENT1HsnpD1OsJos3i8OEjZ+IQo8fElcJKrkn1qo1wYt8eadROVkAEh6LHj/yFa8m+89pQ3mx
s0lpeXcqJaX8TggwOw9fXwvJlMXaXgR9i8VtlA45SG2bUUP7/DO8+MqFPgmfX0UeyW/ZphRee5oP
0yHqZein9OV14jRFDCJ1G3voAmD0LkeANIqf73dQoO4gRANdgCKBFgYQMQtsH/cIEya3CjS0hN1x
GTpK/DKuD6wOhpKQ+mMdZwv0fJfdXdlDC4E34vOynKAgaRhKYHqGSBJfmy1nFaEpr3zk1XeUsFPi
HsHsVhSaQWlfVTyDBN+hPRn4aDpHWZUa4nOn3ibnuOKcxMgDXWKPV9OngW6tAEkye3wFsTMvrqGz
5O/GCKtit1Lf0CL3sNCw+UWDNf6XMGrXx4+5QAV8OLLHor4RkxmKG4IQbPb+804hPdTz+QkVuubU
YlWw9/F+HXhq4tDUzVCbxLcNinskHUd3gefEPIyebScOXL/RUJ5IQEpi7D/pG7o/nPbvePkwsHzr
GLOPtmIDFPNZXLUpl6xUPd0AAyXdX3Hqy/EIXrjmdr6+dkQlk4lbKGxkrfn6LanR5bhVzLy3zTgN
+D2fK2SIb/d4nryKlWfHb7GJ2Y24Jsngb2cPtxSn9gBmxiBoRBSO0PdBXlGmJ7yDofdsYe8Ur1ws
t26SGvxW3w9TxVIsOLdL2HIKUm8/j8KYnaXgwk0f4wW66f2a1crN2Dfj3wyH6YqyKH5inqBxUEI9
hEibpmg7UQRi8EAMbobpMsP0mVNQVZX1nmRB9Ihp9hMLGz1jAnKPYyDM9Fp1TjH5ojosjLARcNc0
WEzvAnu4Gs9jVa0Ur36taambD3BhsjUq1PtQIKamBJX1NTIrj933pf3ehHTIwFK1gIsa20jmrNOe
qTWHCcq4TUy+yb1GUNZp+KsFeSFtUzwHjU6dCkY8MwdL3onBOxJVFOBv0RSdZnvRAs9SJv3s1s6l
q/fcmy/K5xGFMLmu9qA/WjgTo2TW9Z7K5Q7GmAZjm0+JyGGXYbX3J4Owz7qmXpZyhvv5ZmdPTPIk
RkPhqLXMKX9EtliJXgDJEC0FYxLF7R0NH/0zcQ8oXrBMj60cngmTWWmqsDw/QSpRVQN8JilxmE84
PvFluJw2h1tPEeGO3PSVWL1o2N+hgPRE9KIDSt1pfYL9wdiVHUGO7B2RzeRGhjsMiaLwaKZfzd+q
kBKIlb8xBXEaL2VzOIVt88RH1vdKlcMyZFlFH+6gV0ieltYaDrMJtPR25umaE903EszghcqV106I
p0UuAn2etIOdyfiqo6CUh/uJMS8M7B6g59+Hp4I4SwTB9Ogczj1t9DVanXwqZ7M9U83GwDQzZ5mH
H+F/SIFKZ0ZxpfOJ2G5QcmtttY6wbkabSSc3V/3kVOIlz3t1EeMuLsQncF3dDnfL77ySmsBvj1O8
SO0qWNeKwLflqua+vkLv44GhycVLCH4vUYoAyMUEp0wZK+IkQnENKPW8ib4dV3KcKImv9BCTJD9s
FMeIfO0rWoLUfFKCV+QfjC89Kayo2jpL3BLkiLPdrWASegtTqgwk0UXAak7O2AD8Hy1tJF4gJqLW
VCvje8Udiy9LEyDKWuafw/iUj/QB05blTyjmI4+HhtoDf3lOqKrrvt9y6Qt6NBbvJg21KA/8QtrP
dt9m3h/k4Zt8ZRvz+KdZFXOPrrOCOZj4XZiJ8L3xQK4nk5hG6P4HDOopDU5QQhk2dC1ngRVTWV3J
8KWVfEHXfHnMvwYoAox28NChLQjYcF8YrNfeFZKnu2AVMW1M0Hxnw/skGK79pF51YgZnTtcj5b76
6NV9fpCmNX60Ugitm8kP3gDBHig1PnJ5Qf0z8xAruSTNpDHEv2enTIxq2S513bc4VBWfetFwbGy6
g2pbyLz3WoIcJ0wzlsOIxA2ZL0f8G5mie3PSj5W6Ytk5BkEPTotqjUqiQJRpTlmLmT4wR4+50DNL
2ZLqubudxxRRw+K0jOWAx0sB0a46qtuv40jCGM98pTewmI8VO8IeSlDAPCpdb9VPLLKI9NMUKAB+
Ds1HynkEnJ4ul9+tRxfzpcAsR19V2Poy36VLwY9VZ0PxvyKAf7zvme6EojUznhXXWEBOhOol0EXG
PWVUB45nTkmIGEH9UUZsw7qJZM1Vld9ZxdkaWsefsMZr+FI7YEXb/oD2tWfG2eUCewJNjmMFZCWW
itaZ6L8cSwuxEmDKv5krxHgbj0ZZfy+pGjDTxMAPewlFt+W5ilGwxEUVHlXhKnkrPx4yrwQRG2L4
uHkFMTGPsly6V6QhXJmuq8hVkRRpk1KfCWZB7RaE8hCbrxLlhaJ/g952iVat9dhZUWsfOzGGg9BO
J2lubJvUPLXc9HZjgdyScZOUDLCcrN1f9ZNUdvAThce3lkleKZYFev17YCfbXKF0m7JJxbu+/C6j
n5ia+Vs8kmEWmlnII/2/ieRGG4dBY+qH1BU/gLdhXm4hrZGbwE8PV53e4y5mpcG8dAWthHXhChGi
3y45ju5amDtL1Yocr9EWFI83ha1G2zFwnqh3jXLa2UOYuyzfWlzsG9XF/jLUFOOzJGZlli67p7VK
7DunacAqQuqliQ9fgSBi/C2le1Ossc0SutHw3N1ejk+OtJbHvDYNLV0z1OGPKzSAhWoMUjAzLYWe
ZvyRXvKJw5V8ERonlhmnelumjqq2zMJPrvWRmtg0+QV0fF99V/mWM54IQBQtmch3MZ0gyaPhKbY4
LARpU8sDl1J4UTtYUijiNxmvQnuQTWldQlA2T7fZU6CHQvUGYu/DLzigtwVXK31AY/Wtnk0RbNum
tcSURqb/bJNVM+L2W2Zckdsvw9Dwt6XRUFGQSbuIAm+ycssASnN9quLpN1969RFRaH1lmTj1OZvj
f9EG3D0S+pR6LQ7iQKiC9J8q0hNAmGMBN4XZII/f6/6RJE2UOpivu5FQppJYyP4VxqTCU9EHrAX3
XABz+dracSr+fYXfOoOamtqozE7Qq0ZKFdiN/qzfyF8ZKrqe1oOaBT/Gr4NjMTWmxmSPoeymxhL+
KsYyl4RnEae3LXIViHDCv0S6Da9spgp2ObTqpRua3XTLcWtR3olguu0hDAeubD+7Xv+4wTgMWsNy
7XlSY1t0URejeGZ69jc6aoxhjkFOO6y6gSiqapAZWLQLQIURkqRlSrxnD5pkoG/ILhfQS6StD0mB
wcA1eNJ+qD5AbRI1fwTip72ZFSK9yiRzynVAHX55qBWi3U8+oMPZx/8g2GpRPa7p6iVIws7t4DMu
MjMBbNnNgloxSBj67fFhjHkCBT9xYHeIySWTy1Q9hNk9s7QGtGfqzbxKImZjUDA5AcOzc0AzHYXv
XCcptGrN8crgDOF94OhtNz/KNqC4N+5yQKiQdeicqEQZgn++6mHYGh66OMnb8Y4iRWZf99z8ebge
O3CAuAUbOyErY1iXN68jTif9PnPcAL3aRar2RnUhewxd1+meJI0pGA1mJLQ01sL6dpRdggebk1XS
etf2xnL36VpusgR+sKwr5AUa5jc33zesUeIaHijBKf29HEie/Q31w3Kc1MiFvkaBf0oUKkIuWY8c
/e3rxSbgD7kM1pbB3xbFpB9KzJz5/Nfkt0I3YDNwknFVdEa6W3BEy4dFHe7oPihQJqVDqg2aNWdl
qdXj7jAMI91ZdZCjuDSjVGr05AmeS567zt2Eb/J6PcYLTaj8Q6t1Q5NU+Olv4jr2BmSHpiGThane
+twW/VjPSyyE38q0gpgeKvZeZQz5Cs4Em2hb+Jvl06UnovBaiZQm8hX/pNNIBs18zAqEqXpOUcym
Yf9yuza4PYG9V2Zi3eAOar2RCiDxn/+cgYynQR0xziYMKBggQjakgmU31vB/yl8TiENsOK8Tusar
xciU+EiBJu+bzkW3rPf0Zjn4yep6GYCWUm+l1HPf+dX5uXzi2leEL9ae5jmhyQFqnl+F9mX3NXMZ
TlL49rj5mimUPzGQcq4Zh4ggHV35oCGWjx/kEDF9jtz36mz9/+P2GKib/xIS63QTF5bEErcmvC/5
1KWMGZbykUTYO/3gAwAZQzohcpf9J4zVT9GfoJ4I4o2ODhz/TgOyG3ZSjy7z4W8pa9TeaG8SYNns
p4A5ZA7uT4RGLLS6IHVL3LErWjUIciXlNG8fStEJoJUFnFR7K5Zn5auCKMBzMyO/HI2QR7Xtc7l9
cZ/eAWFIbIwFOhs4pwqgBms0Hz2oeiqiylfcEOjaUmQd4KeAFoOSiE2EIBKxNocS/HcG9xYO3MBg
Odkp6fBV2YVCSEOPpSksmYmAeFqmTx0o83KtEa0FZHMPIfCfBr+arb1rkuLO1BnLqYpyGxqDiNld
8zv0QYS0+uldFxgi68kyzURtpa8FUR6v0Qc2yHE6NEqOsimk8VZzVcERWtPwcC5ymCVuW3I7ZN9A
NuejY0ANP4swiyo74tgV3VrahsFYAsRIAam0vScFAJJtTZjcsQ+px1RP7jq//uedym+8pog5V8tH
JntMOzaSDaW92NjLJAUcwTN1lSJjwXxHpMbwpNax41BmUv3JJMeMJmWGywJ3BjLALdXhg3qRt37G
5K50LL+l7cAz+hRzjHmngy2A1wKFJnOenp914BLwNVRmOKWPc6s/njXXalfF4MXfheCtY/03YiVZ
POpiXDblNgZGxBUJlBPUUc/6mTiQOmkitu3bATHKX1OrMfPD39U3bqERR9QvvKKQkKFIU4JrLC2s
ifWZcXFTnFFeTCslrHn/7Ul8ko0g69RTCGkiY/sQ8eVzDUfveLgUjkzVeG9IHMAA2LL9mgdYAYyp
i2vxUrA2egWubv0OnQZKTbFnjfwTQKo/s1rvb1vxD7K6HqT/s4cGeC946OQnMp4u/ESabpxBt3UY
5EQ5nD87ljYZNTnK+Cuhm26RM0K/poacC4fR+ADJyejWYFRGuiZDMgvcw21IwxEZltxiccEartmq
3ijcU5JE5SjuxRuc2H6n0sPs8JGclom9t1fxOK/go8EWaIpoRl5cxFMgZ/Scu1/FE0c0NlZcy48O
AZ8KRsWrACft6JjF/594l0hO341HHW4HFkyo6rfwvQMe5XgNsn98DOI7rNe3DyLLkfnPn+7x9gge
MiVRYifwv4xEOyG9VQut9VsPwLWDh9txFvH7nb6TnqGZWwe+BkfWBJNQewMtUAT1GuyzcsLd8P5P
GLf4s/HkeBcDXHNnQng5niNtwBBdEbSbTYtTljR4XhKMafxErXE+fUOdoqFFDRU28fmkHNEpxjqd
aoFQnit2aSK4O/or8m7QpExAdZT2Zj8yw1nDMamFKXpDnhx+yfXj4GHg3BBdzyMuGZnbgI3RQvmT
VITU1rVqLIwGbhwmWn4J7/jPVTK8tiE8eixuT4o9ZXnZCYECZTfUpvbbTqcQeeL23VZJqzN24JWq
Wc3826ZC6fP+JFUR1CwHW1hb6mDniSC1BK/SWBU/xRWw9RH0oXulstBQqZoQbcxKcsTubapEPnRi
mv6hbcmVQz5l8AR3yu/rbalKgpTHimy82nR1wnOkA077hCdkd+1m2zjeg9f2/seckGsouKGTyIZA
5Wdy445hwe08oyWmmP3N4M0U49SMv9TpnA+b1C7piJqMS/rBcFiabZsxa2/4fN0No/rkw9gBcswC
192Pfa3fFs57CByI2ZPfrOpyyeae6vJajlMHVRbLGmTaQE/Ou3Bq/oPFSj5XcmHGACRvj/6r73Hk
ZR57djpGZ8t7RlrUhmcm7Uaa0R3jVssi6xrbDbfHAa3PM+wnJ1sob+FApgr59i+K16KjdWfBQboA
foGcvyksW4vZy5hKnRXlJsljD4ny0Y1kSDM3+amF3gMKXLI6lbD6C5Dj2p2wMuORODOZmUWS1hMe
K6HoUmWNpkPXfNeyzKqVFmfQNt5uI5IBvcJ9KLkPsRpxXNtjWn0rEoMH/j6CFNWDHkML5ibbwa34
+0DmZZQd0+MoEgkjRZKp5NeikmUBGzbmdQjOa2ZYfDlKmIO1ovrh2DF/Qr6qzwy4N4F/s5dlAgsP
0hMm8N0HZ2FkwIQNRigW9UkQlr1X39rgqHIT0yjATWSfW9tHQPBl8d9hg7xwByeyZ6pncEfTFuZQ
ypsJrRMm3eQ9pfDeG0xg1Pq0hqOjWvpmdF1jPF6XyXHz8+XWCzvcTE3MLHAbazmLva8gUw9xwGG5
eKiAL9hveaJkADvOoiC0+fnCkf7bhh2nxklyeNU2Njgegs9YTcL8BbCBwnciaxK47PboBi4Z9Gde
rm2WMXElIq8tIPuUI4MIuoWIQ80M2G663vCYf2jAOTwK6V1m8kt3R2Pl6dQruSP4+b/GD6BNjV1j
8g54He79vmzyJIZK7gUAdh6ssV9gFp1Vm9MCTCUWx5KtFVrwPDXBtSNijKNWYmen5MRKErtyUdVs
bPO9T9El0vDT3FeZGtiPkPMcpgr7Hhh2S363yxCU53/Df7++I1E14METE630MbSBmeBYfbCADkTU
7i1NcEsVZN3+n4aeb0FWq0JCVVhWyENPe74NwJkQouW9aSLitQLwuAF3iccOYFSCU/j219KhYneX
0pbjtqpjkdIM8Fe4oJzmxymvTbvxVbpZwvKUyWx7fKMWoU5AH2FO1dMb2dZY0rYVvBkxSuUdqaSB
JRrZKtHX9tVxaG+o+qZdcc/X1A6vXNewZgHwE/lx+UOHZdjaIIPBXtT9FvUcBOygKw3ZjwZY/7To
4DKwqOSkHGj5WmRGeoExgigI32gXjqkGMUsBprOjtZkIBSk0wJxIciwx4zz7Wr/jTMT5Am7Pmmax
an2Gnv9HYoqYVxnumogLhsJKYRS4JEujlUel0FOcuEGS740y0VMEmrL3N5ki5NugstP3vWt5bgwu
cxN/A2X/+LMxezgG31yr/R1gr6I5rIrWmg9OtSEHJLgZORAvUCJnTcNcZ/y2espMXwSyfmjB8SJ/
b4qmdO2v5ts8BinoAln5OvV9ISLZJ7RqDxfr11JPR6YjNGW2HMv0FFrLYjL3AJBBgyuqINUMAfFh
PY7v2gvBpSCeJZPo/BfBMO31mF8oLEAkvAC8Ho3iIKeblUSrg2DTr2SwU7o7sxcMwF01mkZRBfoi
DK8CNsqwz54l0WTzTvjI11KBY4xa3gLa0oafZLZeCWczXgmDALTv/v9mWbTW/tFb8nCN45CrJvPW
9sHA4OobmaSAY4LWbeyKWa1J81NHvJFh2R5BjVqeCGaHmB6sj8VPjrcPBJ5VzIAG19t7kvAAz0OD
vlJydAKGegHpKFK0d1bnYsGt4meaHn434w+cIBvqdGO+D1MAx0DMIUBKcBnbF0oTSGKjT5DSsycJ
Cf7gE7FhRkSUOJHRZT2Nr+/SHvfZz5dHpnxUvoSfCDEsXhLanXLXfrpQc7/VdJAYj/JUFizUw124
PhJXSRYwP19owiCRakMjNGDJL5Wh4fr/p2Q+/8qjC4s1u0BIUx4337N2I4HFW6ZnWc3JmSMrbSGh
fhMOQOPJNR/Z/zIfjaIsFxLBDZh2sAh2qKvMG4jWF22sIHG3QUWF1tdBVr4m1ASsiEhoXo9iZXMX
7xL5PlWfAwsfHSZYKuY7prlOBjq46/4YOqxW+3qwCT8KIFsXqdQ4V06smdew0yIGvNL3czpINoqt
3e7LY/JT5bVYMPeEoWaQk03LahPgU3Nc5VdWplaLrrLweLcONjnq8XCKyAW+o5hMV06dx5GqPfcF
CcU3N5o1ouVx02syaD3+o/zScM4O6m+S7oRMcV2i8GLmQ/SFaax12CUpVrh3SKICkgNkZAGHemv4
neDRmROXt0Hc0jmsGR216kP0dX08c9Ez+DTCyqrZ1PZBoUxOZq3G0iEAbzTqvcvpOFPGVQyMAnkF
9X8feOAacFFAUoNz2EambfwaSq4PL9PhZNFJdrQ3We0Xy1rSXOonHd0JAb6ObU4txt1lcQ9T9av4
PJFcGcDDT3jh3EIVDJlVzMWJLlaLpZ1Ef1fkVYkN3GexBDpr/TdbcqX6kuM2a4sY8wHxZngfvwjj
EJDjWW8TFoA5yJNPrl7TooQibdCMzNa6LY4DMN3sWRWcbfDYrAbsqrFnw8IPVZv+Fu0x5S12SxO/
rOijE0YWIZ1ZbdUfVMVjGI/jcX65+HLaTXrjY6sDIjozwlHvX6BWcawxPxKqvSDLGpy9DGOdIE0m
eydJtMarj04vxDoT41vVyP2iaW5VTSpR8WepFHYXvEbtqubVb/8N/vTUbOreBD4ageeO6pGKTtn2
W9LkdvLIIDv7JM1RazPHOPOVw1wG/ghg+agFkVIHyIYO86TXmlLp0xvwW6QRFAixyNivQJTNrvh+
Zu5jOSmmr2NlvCA4N4Ru6EU/S3JsgUyha9bFeRHxQuufOM6LgOdAflfn0bHxOjzNYikh/pAB0xP+
ObOUTgxZD5GeR/4dmvYbYk15Yv9wgaqKvrhnX8chJ6Z8MKS62FFymstE9XvP4yrfieKjEQIj3NLB
sVHgphIj5DomYD9mEObOOMDSY/tkjVdJONQjnCPRk2fMIYGF50TPyApNQEvSrx0/1lPKOppOXvjX
Cd57LzJrZtdd4QNxBwIgGIeSVxSqafCwLhMQddLfWltDK2ISUHbTcAQ2X4s5NGKv4Mphv69YIqXD
JhdcLuyd1hi3EDuHzypFuhhHZkCf35wk3QK6DMSqQIUrB8I2IL1dcfjokLUe6S7VJ2jYV1wA9lOz
yJcT2to3AZM0UdBmTx+qpINUoHEAkc6Ewu+Bqnr3DIeQUOjkqAq0iJNdOHx592Azev9XuX9s86P6
+iF6cXwdEqdLVZwppRSlk+uxyj8fXpJ4A3z/+Qb1YZ+PZm4huCqU5ilMkjNZd4kGqpSFZ4ar8yg4
gmaJg9hVWj9dLGT3IMsOx6rk9ho6+Dy/ZAULRIIp/aGgYE4dXJJg2mbpM40THva8vZxPMdG0BxWG
lFUHpN6WX9G3QW+7W3X6XC55oOKBBzhKjz/r7wHnSFDpyIHnYScNa2j05JrjtqProxoEtUJN//uY
VhD1k4TEWdDbcBEUh01qw072RvKG7MbQqWMojGb0f16PDiPlcVz9uLGE3vx+L7Gqrhhlu0Si++it
1O5uMRJFfBPzzq6pb/yq7N2tLAr5q+ykLtwI6F8vjpRByhiOzW+EzhoD+UXuqQd+pA6A3p1jVP4m
ptle3kvOIlfzRFw9bKR/wyb6whgIqs5Liy+aKu+dyun5itzG9emKsT18eev60HPwrzU7BNP8DD8/
vjYFiLqMngqEbR+fTzNZUf1ffAbZO/3lDJRvcJ1x/UeegmC4G60WsuqCP5daPPgwPTkXzOxtqbtK
FkdzQN4Sf4ftaB3NQDl9tsB/+4SVxE9ieqsGs9wze+jXktKoDD0ZVkNDqB22RrEDsz3446iSCgyo
cSx8hxbmzNemtDp8VDTyI+N9Ph5AehFCpiLJ4Q4sFel9wUCji0t2g4HE6ieyGldT90a0gRoCpfEc
uMByB9I2bBTfrEuHUY9nAiW9qVtCy5MTBLX5WO6wYcBlhcjkTod1nFDRRqnxELK/A/ou1BQ/6lBc
H9zxcIvbq7/JisdYmsqGX32OqWAFdvE+7McI9zaeZ1Iec2H1ySOPMpkp1P7wlBpoau75waYZkCKK
XG/7hZCEL9MbMaJaceY3t9wM68MnocR/Bg/oN5I4SSEk77oUeJd+DF3V6tDGFZI+QAG9J+akn0pO
Zarcw7QtpR93uXi+WZDWvbIPsz24OjmrCgyKaK2WASOyPJ/KSYLb1UJQ91j9LP941Oy8+gDcHoEx
15XqQDKtF8W3vfh1QZPq7J9cMUjFaf+PC4BvfPvHWJlh7G5vxSals/qRZOGjHwH1Lr/duj0dv0hC
UXfqD1kA7pDMguc6tXpjIsOcwXn9kgP1mlLNkOU/CPNUT2O0r/RYHux7CHhHLcFMsGiAEvDWmWkH
mlD9P1kPbtg5rtoTse+Caip7OBoquZU1kL9imXCb1npGbqwoTv5kVwMQwe6LjKpA/DWaWO/Yt7M1
VMnGIzaVeaWPrkGJwuaXNCwFMbQSbcK53hUlIhSGMwhJ0g4XoWpV1D+n/3z26jLUzLF43BDORB1F
T5uLMTQtLJU4ysKHw8OT9gMyQQxAVE+U7H1KVg8pA6wDeepyukXHtJYjOksXHVVNWbWIVKbMxSsZ
e1oXaK4eyId7bzD1h3jbKZ4TPObqAh84wltRh3G8uK612m3gUpFchO3f1NFTTuSBj5M1tuQfm9Fu
/wiTOm0VaAf3/7yibzp/WXQRTJPevm8VsTPHupHBm0fn9Nf2j/7Cl6457kI1/pfQ61OnJH70VCYV
IgqM2LR1nQoov31VuJBPyNK8CHaPJQe3M6RkooHg32k0aeNB1lUXLLqve1DZntnGVMkc+CegtFNq
UitM2znsaavdqjMaVl8222OicRMYYD8tP7xEytVm8eE60Uyi+D6MHhPt4fdYg6fm7EfERCW4obn4
rOoMHofLVsQMNe03XhYza/veGwFoabgM/rEtuyj8gMM1PsvjhOENKSxjfoLs18n9OfNOQCi3hxDC
09yG9kqGlZaB9FaGwcdcwhLq2faZGvt1qxZa4+gG8qv+WCXgc6UEG1rwOAgzikGx8xH5iRCAZhVo
V9PPf0Jdzp4mQHCkdWb5dXc3B513MnpqcLepst3LWzktjkNVWHWBS8Plh42BxdbUq/Uw/tgmi8Z8
ELZAb+NAcpMStQwZNIEeKhOFBg1Rikxu38WGKiWW9Z09YfB2/8DrEQjhQPYbkU937oP1KGb0VVI0
plavBLhswdmesvKhJRmaGidb+umd14cEKlg0ynKg3yqvWjI+OeGQGa5Hq7b4gB53EEEBqV1e9Arc
cJdYyDkxTWw0THaeU5lq/ZnUlVhvNLuT16WRR5Y7/MVM30XggHxl+TKTUoy8NlKc1sRL9jTltb17
noRpVa38H5Vjvz05TBRTfkWhgSChwaR4Joy32fyOEn/o749VftAluvGpkPty76ah7pTF3g7odx7y
eZ8IQPr66ozt0yPdIfsKqucS8BwOLfkguYkBuKjHH2c0N7pME8nPON+X0UxNxCk3bVHEKumC+ykj
g7tMsiTSTNQn1Q0iEATPMGKNFS4WMtHmqzanPehUS4nUIhKu8aaOmT3O3q9hnb/AV89yasDks0I/
e/fp8B79UpXyqNIvNNPApL0ukSsvsiaiodWCoT6Pm2CNsPgzcNYKY+kaOFGc8sG8ew91jdXz5zpo
SXCtAQdHv1Q7AF4ZT2OCcoyinqstcPTQ4H/JKJ6T+fZhXYUnjdHGHV8F2ez+oxDS1rKhYbztdu0M
Q6lXN+lKnvbgL/cR+v5hpSuGLnhdDVmpxuWBQFGVaaxSVEWCM4aaN6WEdQ1DcDH9jpxyIKueF6IS
fTQuN/W/DVHtzjZZ9HdKrjxeVw8IhOD/oOKHeCbKTz7RvnihXkcJviFoZlsuQpjlfEsxsomO8c8K
eKxC0LOSJwwMTuBp/95qnEvj8nfT7pPHdAW5lg3OORoLsRxUsWH4ASeK2mnD3pKwVWKGG2F0xwCc
CszcIXP01UaiEDW75Ol16WtKpTarG1fO0xKlq1SPAwOfaJ/6SebuB1iFW2WPJmTq/5BoTSjyBv5+
zpL6ZWxDD48kB/3BxM8QJUvHXZdO7u80JktFsdbIsKh6Q4STwS//xkC69Ec+tAEUCUJgBvWL5MCu
fhUbTlONoPnaQNowB8KFLDvCOaLYF5x+4APw+bYD9JrXj2OFTLeuMMYS6CXfxz0uWqolBHI2C9/T
BqKcKaen4Tf5EFNc346uAToF8VwSfl+629s4u17Um33+jHjfzNyrtAuLKbdHuaEVSn/OJ3LkC0dq
Bt4oj6zJJpIgqTwA58u8/oCoNChWEihfkJKIICpAdh+4FjGsshtcGea/rPH6Src4Ci0JC/Q++/1L
UfMmDXL8kSnKgGh4dp5mW+NJ90LmuZyJ7TGfKFfHfrTBObB43TaS91JAxUz+xDBrpsQnTQ91GYQF
EeqF+jY4uhzt2MkNpG4rFAyPnuZjx/zXB+MGHkoE9sr6q20H9jdA7aNyw312WPNYncgyHwX6RM91
e5z6LkzqwEBQuT5A1zrDqXcc2oR5l+49q7m1+w7f6G+Fpp1r2KSmXvkTbn3tLM3h1ExRhi+PcAre
sIq1ayIuKnSCuz663++kfZ66FBP0K3iQXklDf2CrKPFgkIhD+eaFbDOj7GcomFR6UGp/OXu7SDqq
7F6dYfgkSXHqsME+3gWnxhlF09Y/jIju9aTmT0FyDBFdJfZ0TtsUZVGxpYGi1Y/kDXu4CCv1Z3HX
P6lKZ+BWgdW2pON+LKGfjiIUEnj5kDXrkeTRJuGxMeit1pCfYmuQkMFHpweUgvhe5KodMAfmJmsS
KNm7LqSaw9hbyDvApe7DeDnfWXHCM32/HO5J2cnILmzTdMQN4IKOMSayZpcdaQyVyVl/uNSOygHa
JZQuETycEFu5PBMwtR24vNK9fieQ75bfIWCaFZD31ESWJTBGCbsw6xJ1KfW7lyTCNE+W77G5xU1t
O8iXzp+eAXvEsVcsZdwlZcMDonoXHu+kXrmMCT2Auz2njr8qq/BVdyzNEFBQquDZGqhmIKJv2+bp
sNMp4mugxgXSAKqFzJyLmL0Hko8omb6PVoVNpF3hTMFeNi3gb97hNlwbQ/863KBWiZSP/OEjF+7v
3Ex7B+PXasEWEnsE2Ykm9lgo73PE8LdfjBDwJaGzk7i7uBd82pNsvTQ0xnceT+FD3Plb+Biw1XdP
GxsHqEPHYCf/SDKbOCvHQYcCmLB/4B8cUSgZrmH7q+1mxRACIya5+Lotthbs70HBMRdV/imxQKtz
hIF3+3MhFlmrfFKtv58+Gbc7j2IIKA0/MOaPciLcqPXUZ7i8fxVGrdnbLuPSpZeO7ssRFVwgJYOU
mM5hYyXGsbrWgwvxOuosNKjqYfSnF4qwRZoFxXhzMiSIfzajBa71JabFVKufyyE4Znt3nSHIkZPm
1IAfHIM51MiW4kKq1+KtLcGiDBU1JvppyZAHXwQHn/08V7qqow6CKtpk8EQey1IB/VV9nlGjDARU
SLaIAlnqPYidhXI1+VzeW/1veB0K0TcEEzIWSgldS37KGWRdkFq6x5N48XQwBhWzcT3p+/jtKSF3
Wbr2n4EY27fh2LWMJRXeDzwJR1/RdC+AdoQtBbtEmWSAlE0pGvlIJRJvGiWovOtQ7a7LPq0RjdZu
3bKjsDqAJOLmVKNS1/jsN5YZ5jUnjm6ss3gyDeRA62ECYg8/TYFu+zLB4LjZwkY1t+gP9gTkRTQw
TaxT0CYZs3Re89+6loizJhq8QayktPTQsVQDg9zLNcf0QLy9ejggAcK1Pp+Be0SRYQ5NOIJjboK+
AMNzKSqWmjkLPrAa4RI9K4u99HS3InEPjo8zO3E8mWRtuxRs/WAuedkOQyhjy3P0n93/Cj8lzmZo
7wT1+m6Vl5GMsahfLFLdKxqaQJSmOmP1Q2Xl1WuqpuHBjwPJjv/PDjyJo4crFax1tRKra+Xyd/mS
loPGcsupt5HrTVdoqnM0siyUKMrcxY1doZK1ZFGn05qfn7fQQbrzlRW4dNASclwKQuRhgB+wnJ8S
roU1D4kN/Ztf00MfSkcVbnyZ2clzGE3gTZThyOvZBAcjHBJ9eYrnv94RxSuv7WT511lTWRn8Unwc
5CTFlbNh3Z5X6WrXL2AQ0dZF03XfAtD4cpxBH9ZElRfxLuF6aV5jmnhXZHg2uNpOTYSDx/iuW4i/
pYz3cOigrk5OOnkiaCFTVvHo6CDhALZKjI3fh30sC1rHLFvo9bY4YQwwAfliy4a/twzYDCqPcTti
M/znmfs3CR08Yy/5LFdATGzyoROh+6n0zXASzJNa8iUWmlJN4iHNGqpImVteIkeP1RR5P8SjawC9
HDtgVDQ+D1DJa+DeUdtrcSLae+dUzOZWjNmosZXMtq9eMkNxfSGaWYEgaXd9278e67KM1OsfSdVE
WyN1VBBFkbXC5gl70gmwO5patYcmfM5eGOZ3A51oPOPJYpVmfO3b9owCGO5XXs5/0P36IM9l8jPZ
LMxEzGUROxafSlZgb7fa7foWH3MTFJcZwnZthIoSYuvn2QTm2rK2CETIe+hi0TAo3/bjogm+eHmW
2PpbNhqA4rMHvz/45t2swyXwQAsSzJgl5fo4A7CLERrVz2ekv1jwOookss8H+lfF44I7KCreLswR
D6QhdX08O+UU/Ce6Hac6YQrUWjQTI4lBEiMqLmhsjjKIfKsHTXo949wqoPWNV6Tc0NtitFa13bw8
b2vC4+c6mQfssXuxUEFndEpSIFZj0CWeuPLzgEGcP6LgSDVEOUWOG/Uts6luBREeF4GUVZZ92RXl
Il9cDM5MPT4Q7pBBGG+1RKrylqrTc9o+AqsIDERNraiDZ5Jfll5h19VK2WmSeDzU/nqC/V/OEOXR
T2Gaxy8vlPMB2bca2WBLd1W3abKD2DAN4zeeEoTE+jGRdkPbqn2PhHr179TEfXgL4S2Wkv0y9ibm
3UJFpXWDis4vjdj/WQGOZz8NIclWoeVUQYpKfxE3HLelkI+3Apkrb0sW22am4HyC3MF4bDp8v3de
nd30wJjXf2WuxO2EMPSsMG0jqHytNlzcXcoeRsOa8U+hkyuPdIjzWQUe0OUECr/ogSu5mYAYdx/m
zrrUlYdEM5EKqO0cOyD4ve/bjFLNApKtZOt8E78PFLrhf+uyuJXpExB09pIsCtBa76djPkOGEQID
OGZvBnviAVqJ19uZmxMUsNnXH8h1K/hAXBgvHHzUc9wVlwO6fUALABXzelpOpavSNs9OzD5YMDiu
uL4UFKfG5lJu8v9+t41vdJBO9IHznU7ILYRI7cwMyLT3CuftACFnKn7Hg/oRj5CkQngSt+GcHT9f
kSXgC//omFfRMgRGui3qaRNDyPjTp2knilTI6WLHniezBJ2xOF78IOn5W8REOQkTehP5HkjtE/6k
xLgObheJ2Z6YeXyeiimdvePp7VRQlkDbycXPzUAbB+CWSL/vqrrG9luTt52mlxiIaOVrTH+Zp/A7
lnPIu2ZRbsm25DdAssqhHjYI5S+NbUNjSWpBX/wchmygCWj7NSKSYURwx6RO9kBvIHcQPm0oG2NS
p+ZRxzfLHpgh5euNXbm+0gQMNQzygVWWYFS9U1t5VCMwPsSJtlmyNIhYwSmPtkww84Lj7L5CPtSh
ZqogNJP3RK8L/oQ98Va6h0O0uMQrZvkM6um1oFnYDnVQdWlGitdSGPJo2gKtDPQMa0HiiSOLcp4h
qrLSxRqN0KgxA4MNq6FO1QlQ/P4jum8oF2hF0oUu8/UNUM3Vc2p6FJS//SDDO3rCsqPhN9LtyhWu
wG7LChb2awBZaCeAWrvO2NpyyaamLqrCOtwqhfChdar+L53ieQmJsP6Pi6hoYtM91fQnGxWknia9
b+LQnGTfHLocA9YNU40aAI7W7AFqUSc7H2811daEVpstgqDnoR/Lwve2y1Z1b7h/mTSaxXoPdOtt
WEwARfKtP5LXsKRm9s00UQSCZfK5LjziXMMZKWl0vG5Y369Ce6rqp/eRqLYK61hiOTdmggOoYXSw
a45VGS94oNQEfkuyGbrJC9xuowHSoWeI44OB9JMTaRwKMLlaAhVIh/YbqSsPhanSyuFs0Iq0DdcT
daZMvdDG/kzh2bQc2n99OTIzMVHQL3+JVimG6ru/Y4VtGdNjRJEVmdMnkqPR5e/x+DdsZMaSBMqP
l5Bv0HhGw3lvdX/F/65XD5H4aWAbsVJOSrFEQdRe8RareqstrbRhWGRA490ptsGN+1F1UrAaTpJu
0L1t/a6v8eK5bz1pvBZfP9hQATYI90inrT3tLiXb4byeFbRGmZEZmSA9JUQQxtAnIwswLUOhpEge
wzigiiP773UPy/GX088bidopBigAgRzFRtNhW9k32mw4pCh5X3ufCg2+2z40s/Vnoa5gEMUNgPjF
6sjTQXRqLivW1FB8aA4jh/YxAUVDp6d3XC20U7h6RhdkMRuyn26cLt5qFooJY1brUbuLOru8ja3Y
DLSGAJH4DNIxY4yQgfaf3FBigPSXQ/4ggv04VCvsvrqu+KLB/RG8Mz9/0nTlxOnghZR6JxxFvrAE
TbqJ1/PE4U1ghwEPuRRkmjfZ2MCh0aPyb2e0jjny2h9OQIcvEVelkqwFVLUd35GQ/0tu1rU3K8YK
bwpzXVQyqXSQFrwunWsHcN+yCNdBom+AUYLLYJNbXCuCqVysGiPjXcr84qeyOObCP2+bfDGxCriZ
U7pk1YVHNTdHl7ulmIu7AauEIAeJQa5uNrxzgv5925UyGn8VHQrjmY7YupsniTvAz9hyOJE4JxzN
ZGiOIvQ4x7gMXVEGxAyOFTCz5GIxmQxdTbcXn+px3GW8iU+CfwUQ05cB+Ai8d1QbKxq8AKlRX7vU
i2XecD5A5xl7fRjtpFJyIWWfEHvSr8uYm6IMuRpxHYXoYvt/bpT9iUfEm50j2t0YyvVEpAw8ZBm0
U5C+g7aaEQXOsrhenI88uBsvpF3KRfBefXtaMhBori7i+goU0hFEgWpKXucRm43PLf6XfRUJ08aW
+5MLt7rDiDClm7sumLQ51zLdOO3kfEHeSp2D4uziJ+vFiuWOyTFvUz/teiQ6MqInD0wmHfF5cRr0
DguTbLzGDsUbtoEK8sc1hWVZ6K4pmMBayxO8Bp3ZtyQHz2zh0ndQ5vx55KUkfW2Puad58GC2sLO3
EBD/aAIO17Vs2wWlzXc5hiL3JqGvmYX6lclskBto2eH9dv7meGIbZ2rhokdGR4HaxZ/rd25hwDRO
0TvYlRBzjzqTB5GU3CzC9jh6fRY80PEj1kQmAY7JdMuIvzZcM1/Rndi3Gs9jIhsX5gYsTqBUEUWD
fNNVD77WCz8vXbU8Ln/E+rlpVrBRSuxO2zvfcOIPVY+tGO75HbPkl5i1DhFYxL9Meejxr7XXjmOT
o+Sr+BO1jlY6gsRC1MLbITd8vXO+m4BRRf4SuepXhbxQhEW6GKgDfLn3esrBvMGnIMIKtEutSliW
HwcjUWnXQ388KzSEpK8/zpEb0sM622Wmw4uFQJ0KR+DzT9SvvQ4RzE9pWZ66htdqjpaLosQddghO
CSSMJnfMjNEwSzgB9tGEQf/FsZavVKqDDu/USHV79lFmFAxtHeZoHM5DSw1ghF2lcscm4Kk47j1k
oalev8c3sBR/e47v2VKqtaNItEPez0avnbrK8HzHfZ4oeaTnQgl1I+12hPAc5kmZnLmu/wsfCflJ
9BGWs0Cz2Ao79XO8Ks45TdG94tUAa4An6UCzz5o3azKS3VUzcYilQcljWtBcRvi4NSO8lNvm6MoS
TIRYesLEgqIkmJnttQLbUArTuFlRWkR2PU3lqk7XPxwao3FXnSQrVI3ay0zNG9b5+Aa79uqkrbWM
aMyvQqfmtzZMNbfQGFQdHzApg3EytghdBZr9uwf1laJinGgjJLXSgUV+JIAJtpQKihdTuwB8shQe
76JS92VCv0nkewr/s3tjDvitsLLcOaLpD/ky8uvAE7LE5+fP6VG9+2De1JvDfEketefEQj1uoeWo
t2Z6jjr6WlDB/qpd2Y5QUjl2AIp+9U1WklQp35qW1XEIHU+8kboer0lmaiiTXTlPeRHM5GgOtzQO
5ENOGq4X/mG+aYJ+1X9x+MGEZn+7PzvAMQfi7u8+mM9+zxJA2CO8SUG7IQg0++4ib4lk3Nlxm+QN
pODdrZ/nmIC1AEYwO/x5X5CGK/mrDSbxe0ptjwUh1v4I9cAnVO9x1PH+9xmi8OsYtE2VLD/aDJGS
DoPcRA3ylYFrc/WNprB0mLJUtfnuAvvl2MytC0Lt9LHrgBESYw3zZ+eHXjAQE9nu8iehhuMPQ1SO
4STO0JiRZhHu+6ZdvXaYcgODMzSRQHU7Z9YsLIkepbwVSd1hycfaDipDR3sWGgjTn6+w37NUiECy
8oMWG+I+Ci5xCtHLae40lTebE7P8CCIi5Io1afzmNhjBnhnK3Fm9CBnAdkVAanAwbFwlH32Y94eh
LopSRAzCsTaxFSFhXmf6pzDJqHGAY0VKld8qHJepqq4PCcdvRCqF3wMvpjmKzrok6JYDKD/LFdSu
bOMmWylFXyxD6+wCaVg8RTLkA6N2jx2a8zuIGSuEdzPTuPrsyIBbvOzbs6ExOm/P5SNxSreau4Tu
tTsI30G3rf9Gm47+7Dgy2xXVc+4u7dsQKGEcdagNaUwHBgg2NlPNskp78D9dBUnDEUwZiQzEfU/P
56AoCU5h5wM5nwHKz/RtJbaFpkQUdYbdoekqrE84sfXU7a6JbWV9PbncQDrR99Hb2SZ8yDNdbjKC
Dm+Iv3q3VNC5f3oQt75HBb3oIokj2ycq5qdlz+tN9k7D+IEuXLNLr056yUAu6MnkwpeSW8tBSzRZ
TxsWHbw4Nhe6S+y5WAaT2qwIi3UrJALTLkiOlDKJ0/tIiN8Uhjkbt+P2WyI7RA/gvlcYGKL9KRsU
zzUl1g1SnKuhV/rNjgvqt9rY1etT51ZLEJGTWLSGAihNeTwYtLndAJfhzsovaFSSVXfvm3xl1WlD
DXoG84zKL0+UQfOb16sQ2p9t08QeFeONJukbVpgSYg+kcCZXAH88SyJMat1thAaw9lbIk6IS9xPp
i84OkkMomSSCM8o0UIa19ypukNM/N3x1iQHqRsYX28c9Cr5PiZdo9Z8vbd6StMZ8ZEYy/Q0cTIJA
VAkux0ovRqqJk5QIWsKcAwG4YKM+mf4HSkT6590gCo3OiW8qXIgkUW2aYWwxHIlJY2FSA4v0U4Y5
kuUcG7PgZ417uLuNMsJyMeq9zQYVA+wz9bD3lCI++6ZUSUBkZwdi8TzVmO67nqsj3S1bunafhQzc
I8Ubtvh+04/CkAEv20BIDRGaG1dH7cxCSkRlXqvfHrqya3cf/FTXFxDco4T7feowpnCTq8jf/dPU
zPIvpeN0KcJAmcMFWvJmLlmnV62t0bavhW7+30j0WB0ZXwCuja8CiYhPDZy98gNuejDgbaBcYYxI
HP6GX+U67DBZl9pOdzWQHAUSu2IEUDmKP6FW38WqaeOWNCmuZZeYOL2khMgu6QzOL1XNwFU+8X4C
4XqjO7LTVjeJJxBHuD4ysV4rMv3r/WvR8qXXBXKLw7W70ixPIZmQSRWLcFkPSomU6AoJU03M5CVK
s5xG5b6/Hrepr+GqQff7YLuBcSb2r2kw59EIq0zrMKiAOC51L7KZkfQ2lH3IGF1UWr41dMKo30/B
RZ8GIJVQChNDVxcg3zK2ILcCe5jlILWQVbxaki3Yy/REaEhiwNvThf+hULl1W13d52HzYhGSpU/m
DOxj/Ul9rjbzIvfHc7cnX3HYCD0OakqmaWd4tXcuNjoqy0VtiNj3mXBrbrGKMDuC8NPzYRRoM93Q
KD0xjI5aVt38kr39Ztf2nEoJT80/drzD19mZ4VsM3uPlNbCEZacoP+ITIpInZdxT65Zdj7ZOSec7
PMA5WPAEC8mHf1Q83u85Tzx36pZ55f+CGKUdyIXgB/hDhZ7SnPFyFmPDWD7UZ4sRFzUE3emNjb1N
TRiX6SbBPt4zEq27oC0mGLI5PkToxjO3QGStn04u6ys6RQyAYOOOcOUlOUXZamdG6wezgTFZkp6Z
+MVPrJ+OyPEZ3rm/a6FCSjNIPaGfJtmOaQbj3v1UWOQw98nNi+uKkUX7+TP7y9/wi/Kr1pb9sSVv
HL09nSllZbiVeG9lu9z+dUL3l2z1lJdU14Tq1kpZuACcuYEg1iKlXhjwS8Btws6vWTwZLi96+egE
cxbEqpgKjYM7nUejblYlofoe2uFLnOImy/9kQj5UmpMwXSOc5cjgALMvTHJJ/LnvhLTWsM51qPoC
1xCxhFevcagFGSPLTlfSC6s26jHvMsZ82cVMLe1PX+kqfSRhaF+Fwv/Qhq6pEBbfSvaZ8KI9A0tQ
sRG9IeAPR7eiH7otHXWjy6wTNz59n1ytAhQojdNgFYZT0mcmcG7OKZR5ljXzORcjiiBL5yv5VVzR
ALp3k+D212vN8SnG6kGupHzk2CAvwamUeajTT+5HNpr0T2KC/ObN1YoH9XcGkvMC+5XQrYryqi0V
RK868ZYm2EtRtG0JepaTfI076ANiXqIIgQmnBxUAi00/d1lotn+z/EbPYDAKw4BId7abmRJS482o
/sNcZPrq8culo1eWABmoO+5417coMab7qzS1g3M+S2O+Y8b2om7PVM4ybvu5IBf0peh6+8/zYMG1
8Sw9nH1qErdor70Jq85D6rs7hUHlHUCj9t9A9SQPpbdeMfqR/nQle9nzz4sE7goHg9cf3C1lgV6F
7rMz9aHxJWvjZYdcBEMc31UwV+NBSQmilHAzRRxkcVziws5IKI10oBJSJTfb9Aj+mPl3fTa3fxeI
3+2LD3LZqckbhKohHrZbskdTNWZ/pFzAfZ/7YIwGqMdnQ3+iujCR/NNNmDFEAMhKgIuE8ulf6+kZ
Bqz4J50o5GzF7WM8mW19X1BxOw4AB/EIHnqTfr3zk5Ej3ohDn9/mf3dD5EpmdhJFffrpvfk05GPT
7truc5L2yEUkobYRg8TGx8ytAYzqChz+KjJuQ7PGSHxHNikEBeKancDIjU+M6jQg2gSYtW+beeG0
19uSyGJHWaI27p5KZob2ZEtHNZCJjK3br39kdZ7UL8TjT4yPmE2rTfFt+ehjMJP8CR/x0U04eoLg
rlQIRj1KAVcCkDl2JKzormVWQncJOsyRFqgv4lJhyVeHTiRn2+LJ7YXBwRv+VnH/AXXJyj7Cq4UP
FAyqxv2glEAZlGgHC+A32VP7JTxoFhOp5zDNlP9kpGGJYiYV7uMmX2ikxuCsjshR6s+uKTzc91Ax
DDQoCqHmnpmjggsvTB8Gt1dmIV4CWxSVsHaS0oJpOj32I1+k/zyUEWk4qSarJiZ2oklARSgjGv8T
B6mQYzqONWIRujLOSG9XtSDJA6T5O9GYOMLFrfkf/63frv5ciMTmr8DNsDsHIGorarg1YcE+pheb
hnV4mRxKkKw495ajm1AkZWiGVmGqDfYrZecuAKUBo7ccOyDMfyAMERuGAsId93MeAkeGcws6GMyW
Tm6x6FWmz4Akpyh5QHHY3IuUBffhTy07FQ0iyfCHCnnH/LSBepLvOtQIxTIU5rc8y10QReQEW/wE
ymHbYArRKA6NAQzY+gAp2l9ZB161+Y4s7gII/IMf7Ku0ScLNL0+a6tn0Zaxmh/sG6smmkPPuFJJy
lIU0KM7HZaoRY8sNJQ7GqLovoCJ6t3iboohkYsGWm40FDHFVrU/SlHLZVljfugM/RjA9XdkjGMhg
JFsnjOh2NoGTPJtGmygphh4NWU1lnv0NmGuvaVlzq4HedJeASHZqlaF6ZSm4XhZHOHjgZ9p0gtKb
xZn5tvh07TuypgWgruqR4XRKYQkVePKLYnjGWfCwxcDlIGac/wZdr5C46lheYXItfIh7fzJnb1su
bmnogWUAHKFh0Fq+TAnd19Ze9qFPNO/pzs+VtLa5nfpoZztqllcojh3OiuBgrXjXcFSMVhUeAuMB
flgRPiVR0GNTrxkdcThxBGs3jNxsZMLG68JlCyJKhBPbZsPkGzVJPu7xZDxhJr4ffuRQy84EuoQd
tf5HM0v5D8tuaZ6VvjDmUJnd5RpCT9OcNIT2XY2W416yPGe7jC4Bs2MaLRy5ep6WNz1YUF1g3JVc
YbOt7mM/0fHycdOBAcZy1Qo87fxI2A1AgF7tQIEi0/AH6QrRITzVzkmUT1NLtAeZ0LQoIXRbj98X
5f/MlQD2UrkwetkP3By23xEeN83bOoqGVP/W52XIeU+yX0xcmGQMJpdkf5LJXqg5R4Sk+siqkCxw
K1LflcrIdsQSzO4hC2oZDsOzhecEyaoY4VZT0YtkE9IlNJOQnsbS+jEMut/XoStpQDFcZjJ1x+wP
FU2qvCcGVbG3YJAsN1BLl0Q00calSqP1LAw95B902HRT0QoeXfjvuxnhQRBBUCA11oTvJXCJAbhX
f2VMXKE7ffm/rZRtRYPnxQoV0W4Uu4m8LHBRPMRfjSr+ANyQ6ZMxzYVLiDobnIFvY2uAXWcoYrYy
1IFTKg/UG+jK15Mvy9y39J+mEnq2bgxypgxBjATcO9JVEUf+ahfn/hYU4N+rvSoFx1ctnKXlEI1c
fDwgzcilER/MPFX4qbh27XC2/xftWxDBM1EUx70l1wjn94VV2f6UXHPxgSYGqXXnpMbUsuFFQIe1
xhzpQd+ExJ2jBxlOvQSSVGB+iKmXQOUU+5AfJUMdQ4BnG3Zqnj1lNL7doiH1pQU+0t1qiRJz0IT3
MYHKL2b5ZB3DxsibUoDrXn2BXFN4bj6SU98NuCS8cNIEhTh3c46wi1apdBm6s1xDVRyB3zdYX3Af
HLYbunaubWLn9ZQZ1s54C3Z0yBIu821jfVaVHfl3Ssqvv8eAYPxwWz8wmkmyJjyMJfQ/nYNAwoMB
sTxXJhZNtN6r+MjZWOMXP/sVtZoWP7xpaL4WX+62E2ex0MUahCXR+NiCzUrBQ16SQ4VNZB1AZEqF
5moez3Vwr3qy3l0sFoiQ4qG9nEEef2kynQJR8N3BIEb9YWqwwij+hJ8GuN9bEEEDiCxI+DK5X5fw
vcFltGlPWXDfzi+gis6EwjfeSvyiXGEv8iNRcitIMsKLSuPNoyuq3kNejJaWObjIMeB1NxZuuw0h
Q8XdFwZoRWr5rnJPh3TyL/Q/RgBU7RK86nkPqstuVagyidXFVAz+Z08O94CSKCDkWXnYzidqLEJW
5CsPBc1pNy55qbp0ZqncGgIQMmSTH85sxLICpU44dHJuofHQhFTuMO2Q4TPnXvjki0RQ5FpwTAO/
yED3q3yqMZJcDblCu6gEtMWTse38hE6yVdt6V5CnD2FPNTO0h7WFmuAkuBMvM9ecpl5D5z8Q0SdT
VIQgIeLyBtR78mtoL1Eh0YG2Yu/+C73/gWSlQxaZVGWC23t9eO6Rmrn16efJoxndb5VKodyLwcJF
6fta0qmH3oqECcjKDkmRk9Gcqs2ovysQP8iEr4DGoztjFYcmyJmYMYG3Uyp9M8ceWdROE17X/0Ex
XbwvYl5gTWb8tygqIwSrSd300Mi0QXPVqlYb60Q9siwnjRigog47gH3ucNPrkJm9v3JvgLpDTsxT
FqXHRPfhOv+jL4jPvcoWx6bqsdSu3irFXA8x1N8FhKwdAF4lgYFVM3h2+wbCB1RDV/fLfeUP+MNx
P8qZdmDZPmhFe0V7TquLZA5rOkrHhpLEmfVKwjdrD8cb1KKQWbeZJMDw06HyYt1uQj8JALWhd8HB
9O+rlaGzSgN0OdrjOAYto6BvkVA4bhaj/MVc7jSsDcU8N9sEqMQeDQVvR7KVWibuBCN6QLrWVuRU
BqDWfB0c+S2ki3z+DPykVwvNnr3P0ho5xL7GnlcXC+tG1JV/C/8WUw5lf4j5ID9VOwJiFdob1QfW
XrIOCiKTipKDix11jl3YE0N+Q6DXwTSK1kooz5MyjJq6fQxWL3jRXXJRgR0uFXWRHe53mSz/hmm4
O2164gXYXFztOg1ldTzo8urNw6nF1/dDthaeLyLOOVLiLtju0REuRcN6e2H2hoZoUG9rnVlH4hCE
3TRTbgHaPk0FalfH7bpdEW/OzegD/RoH4nwtinSXMqQ05rwGdVqon0YlTST+8vgtX7HKe6eTFoye
pt4IJVm2dD6VtlJKIiCgmaDcisKkhx9XWZZgLhhi5VU/OtdUYAU1lbZUkZ2L25fC0AXn+0+tYlB8
8yq5wrqUFgbWFh6OohVWiZZVjaMUi24FkcW/+3XtrrHgAPJdnadZqQ6fajhlqIgDaHVD3l2PYYOD
+CYg8kucsllZMOpIpdOV2waETn97iVqa5y7qkq5HdLqgxX0RXDf9pQwmnILi+DHf/SEzIjCaxplA
ypGkpIWmH+UdEl/0CB4l2w4fYY735ZAe11MqWq8LQdKc/XPmuRJJcXygWl5DsLfmAccVXY00l5m9
vicAvZq/xzPSkLpZzgfLbuJddM33e8a2igUTw8loJ1td8YK6vciOuYMS2ivx1GpMNZ5kzdE3Cz3+
9NjO0dRjJcHCHoyV8VFeYkhV+5VlWH7RfmW8FFcG7Y7cbE3fQLG0g74A+lka2Yjf7RlpXBXQcItn
fc3cHrreWmSlzetsCPvNofdf9Rx9iZKOnSNongRRqgDozlmrwV8UMk7dNod/ZObYFsHhBKDpp9St
Yj2Cb0A1KQaMm0wSVo9Hh2JpcdARZv5nz3AFacfRAmDMQ8iFHp6JotK28Xrv+zrBns+JFgMdCLQm
B9uVxtVU1jdHJfyxFEM9/l/yE6zLt/7hnLkOGXRkFvVD8OoxLbKtg7/xIrClV7k5Hj+5XgoDXFgy
8rf4nQy2WAHtRRTOcxnejLJapqwz8jAeXJoLmYlvKY8wS2ieQuFEkNOnKTuRIUpaIt5N/77gF+HP
X6TS3Nc9L+XzSkBY6RfcCPewSMTC7N4DOG7VlYj3emuUXJztLYKu4gImWFbNH25T26aEJk0h3OO1
hjdde1i+aUYig/EvKrl+lN2aaJN37TaH2QdJFlQ96YdAQUHTZiAqlv/t2UcbDTcXme0XVs4VRECH
icQBfs1PSxf2DmA2We4lH4kKiAxgq4o0SQwwAPwzAVy6Jak88wt3ZG4C/v6IJJ9JuU0nYDCKT8v+
e2bQ0pnBpsRSDgf/qYAPejUiXgr9N3t9vclx+mGkw5CpblsKKu0S6LLykxzR6i+5B2PQdGg+BLk/
vuz8b+1JnAhzJkCbQ9MZQAp/FpNmKZqjes1TiMRBoSs6+QqZcR4JHXs44ITN1Ouj2S4/Rv4Hbt7l
9n1OEPIMq5NTfx1LB30RZqpIUFoorsGxIesvqtu0CE87dFLNur/xewFX3X3+xZIMzr1SeNc53Bmd
+UjynvYqQVT9DKsoIHnhSvWQelAi70Fhx+ybs4fgxObpcfI3ksWEVCMWeaVArimeYp6Th11FZ2Of
vecRlkpy96MlLnuHLhngjOZlYq3nPNF1gQdfgv9DduWicwY5EtuXZG0qun3BMavyUCHAJyhLHuhm
hinoI1jdXHwvelxFEU4uAYsyQkXwEnUEIM7HIJP4smojP8fsYZ4fYsC6/zeJ95Fw1SAL/C+beoao
4kKyjOte6+FgdsvRO1u0aRTmcfBU2jIwm20N1PUPwzGQrMkAmGAzja+HMSe+Z1fMDXGYzQ540Jmx
yLLiFPE+YnX8dEM3OXGVHANSXHY4e11WML6Lmxw3lUWqddHDNVEQOgSAUt8WQrEah4kIXJVxPyqA
E1CBSxlJeFVHZTdRIayu3w/sAibEJSa6YT41tYx/2ot39Py+Fhe+QHqc/2PnDwtVdzXkMtYC33VD
0qq/ikciKSkrLBfgq54W4ZrQgX2IdXBUwhNs0K/I/AKX6S0yMLntELVo+aVzTAqGzlwMkee2PxOu
JTzW08Jtp0Hr178Lap1X1gIv8UNK4WcFXryCBNQ8K3O6ACMgmt7RLeSyo5dd6XsgWff8UuROTw76
xNH/klaTRS25pinX2hXN7ywkSnoJu6GqwYwWIY2CyLL3X6G83hbjU+iwmMyALQIHFHZc4GP2NGH4
GoBYsDhjvb/fpFg8ygpMMetLDrTfe4b/g3QnfWPFof1HPMW+QIAZAH09EMwPH8oTUdS8pqV4hiHs
fqw+CXxiza6JvAdgNzOvfMQBpi5Zi/ByX/POQgxvf8fpB71rpyVO7NcwnI1461/4/0aHjFlVPYa4
aHElklQv7ppVd+viV1qt+gqlKvI8jihwPvG0BIM14d827b33kxPPrMaABvuwFS7Iy/D8oao/ab5x
hwkPi4OcTEBoxFw1R8AodY1VzThZjzvHDn8nIuydKuJ6hB2Y3ONpaaTlG7YryDoRRD2/bTKptfDN
8cAr0khlMJtHT+zzXc5OUa3CEGbmF3aVi6KcEAd2Qcu3lAH05NJhnW6wqZ2QaabW7w6m+cSs997S
YYQSsOcqIuPHLuaHBp1r1cC8AqMpIl/fv/H+2TFnrU74CWna+ycP5Lz/iMv8a6q7TPZEA01s1a/V
b85rNjprHpVaiaZoYjfm9DpxuCnwHWgg3dFNHV+EG5hQ8VDo4qhaAphDrVePo9LI/8OTUgBN+meu
a6Tmh4FeYfM3iyza11JC+UAojLkLINXbggVSwKjEpPI0uj9iplOiaeBNkwdMNpAI1rMyARHD9lNQ
yRsYpSiaqmw8AbncFtq6nS+xd+gDzhVnkcgmtEU3xntdEt4jxmlugtv5yrvtWga0O2VGaSBqDrq0
Ze1gJHsnXNwVKeYTiCQGJ0aS5tun34+jh5YvU7xkloD3qZD1sQ78QXaWCVVBX9+FbtCdwIgZuCEA
Ss7dFiy+JmqUifgl27tbPSrKKzMO0WDgrqqfpUFrMAsyEdWWSZ1LF7hWdZj2RtLqZ4FBB+EP3bus
yXuaP8IrSeUfGMhd8YMSqgNll4BjPVKQ0MSoJjP6wixQ+5GT/iNgcLMhIQBeHIS51tr1H/v0fU3B
eVNktWKgUOeSxTWA8vZQIIWl/BmYGZqN4tmTo5iEANwsBwkLnwOMKMpsBuP8F9wRtql0spuSb/W+
Zj5HtVrJpulu9lRNK5zyOMcUUTvWrbP7c8kCYc7SxLQJZj2DtR2pkBS+u2Q7eBYXhe9Z9a5HZ7wy
nzHFtTBycmeXdFZeWye4qWNKY29tv8fRmBypx3csm/oRmqthRNNLBYj6Hyd0aB2OTuMH7X62Tdtd
DPjazGdQrGCnttWMK5r944+x4jba5ClJOBcbSUVnpvB7xZMSyjCJEZsyZpJWWxAzibExWOLp2Erp
Pqyhvle1husjg57diQes9eptUcxiP3u/oK/uTsk71kp3peFMwoDVlMnHFaFVsG7CAIN4pq41+tRz
7AJ7m2ljSLSei4QREJku9TPlw7rmwUhO/IfXbRXfz4rHhDeXGdGHh0PuNJsL9bi++pYdjQ/oM40V
WEkzgfJNtoijLVVg2dWWxZkJDft9PJDRp3RQjz12ZPIz3B5pAb1gIsR+y0Nxnb3hp2GLe0TBp7b6
V+80VfqjQTAjdzt6Tw/aX1cOPCXANRZceD9xvydIkGm27pogYLzazva7NePibH9stMemVLCs8kwe
TMbPvuoVeWR3LA4CfZBZfYixZr5tNeBh0cNHo98J1ydtKekXlzUqczjB89JgLtQFT55+5QpLzGaq
MwZ1lINXqjfCtuoyiY2D1Ln+qb02G9p05opFIpvZ33yoLAOGrIsIGbzCbFb5mTv0OLD1MOzNoOB4
7fFNVepF2LZFBdYGb51X5Nivomy3SI0WrBdAaTx9gkkDA2cQ9T9U+K2QR54+1wMNV8Y2nqE6ydLL
MehHa0tLQwl7Rs3zu6lLkwHtgLlfxgiIyr13jt0DxqKaoSjQ7aRo61LfpNEIMcGE7qNJZ9cs8iPe
lJ1kRwHevIkEeJKkA8hjgprDkweAuLuMHv3Zyc5QW5BIbse6/tXzPSmodbaHahztM2U6MLBjkw5G
bbrHeHnsHJTPzJCRFMB7G6f/+EMoEzOOdXr+3b8bPht8mci6IVEaQjNvp9C91/XdPiweC4GnIzSd
ADx3zLEfuOMB0E5bqZNs3DNjx6foWAjYhEa7hH58VMBdCzEz8O8Z9YHuzEk9kr+3QaeEVSvC6TBy
oJgU4kIpNyYL/1kF3kNZIXmOU2eBbrUuGiHxpfUD9VlciMOUhBp395uLnCM5P6vXpN4pWq/7EvXR
e6Hwi9eLV8o4UfpFCbi2TUOz44aHNYUmEX1woj2Zevb3F5X5b1Cjmhi2asuI/GF6ea3ZS0bBnXjp
lo2Szj6z7KjjuXK3XhTUD90u55HX/Jtvo3hewUgyxcHPAhji93pBxVuUB3vysqrKHFQukjdHLfDf
gb73gyJv4CEfrDZG2eJZy92yOP+LbHljqfrtA5UvK7UDesJ3Qhu6tlXgt/kajrAsd8Z7eqxzsD9t
qqd4m7Q/iEP074TVvDepdB2CNgDr06JAnjTuWDt9WlbDLjeG9rRtBiXvSR1DRcWrgLYo1m4MWcmb
bFKRvstGwDuFK7+WAfQO1zoCZnuS9PSy+l/s6t5bbFy0KZ99GvFN3QKAqC6M7KQO4oe6XZgO0uUs
T2VRGSqsFlipb14uovxzWQb0UeJe4LanUUFeo7TSHAFPxvjHHYZd6HT03rsmqlxS+OubKrD+Fp67
vbgnGfyNcHmO6crNvJbKft6QefH05P5W8LpEXno1Y+ku7wsN4eBrCnyUnww2uJZwDPeAksp3tgQ9
da4jPB/nfKnoU+72+i3N7i1vvxyS09yiwqUA3KB6uF7SVOpEmVa9WdxGvd05cvQAaA5jn6+765w1
9T+ovMpVAxLvQ7D3YrN8We6lVOLUkTHhK7ZdDL/8LLYCL+V5pE4a501oa/HDOP2XpYVT9HXFKKJM
iPKQQaIGO7o9d+EUI5eBO/NnN6GCybezrdKofLpu6FSp5OX3f/TXdP2YdS4C2INtnLDMgR1+mHj1
g6FvNUBPUctj7If1DLc+oc65Q8DHOA10WEIdMAD7T71P1NNepLByYvKMNm/fqp1R1aw46hxi2K9J
j0OWsbYURfk1QKB/GfAuTGVLCv/y/Vt7aPgbfP/kB2GxQOCdhiMD5W5bwf3AkSSwHCsraDjE0pJ8
7MsHTgmbqu5jynAIB45O1M2UnIXOJXC809WXkQqV0Ul5+CL1cxGnlg6JdkfkgnqOU+dvnEkMO0jp
+PNxnjWMo8Wc4VTuE+TV2CmO9H3nxUTaAvkkBaxlqhHugsvJVgPyu3PCDUs8r4vtyeT54Rs4CNSY
5Qy7VlmmtchV2ciCstEtxSHLH7swUdGrdmpQFWOBub+dZ8KZGba/8wxYHIJnV6hzrOD2Gkls/+vA
NUrINHBhA+MnctxrifYcGJ6jY9uq+8SuO6Sf4j30THp49FXItzp5c5IzSdDe2KptNm0eqfBTeGKv
QKmEXHHr7yoKO4LRHg/178gmdXC2u8rK52d5SEJW2O98C5TtCs+ZZKkpetbAvsG51BBIJ3SDBqDX
khHJwzW5HahanY6bdBGlBqKWHCMdXYb1ZfoX6hHizUKCpfpcLiufkDICuAyNBt5FA50vDMz1f80d
Prx36qF3/0vTIcfgQesPGOwCIydZIDCUYY5VFHF13k2falpiQZ7m76rWps6Evg/f49GWTjDcS747
iZKLMWFrdVOJzEIBY5AJxFru37RshIJ8YDjnJwQdDpn0kxMFZcx3nYBMOlpufISzrcxiifNdk+oh
B/T8ef4igOx5Oz0UeA4Tc9BPPYBAEtuEodM0IQdI4yXYMxQK4FkDihiZUlYB+rSIlRplN1dt2VU1
hPutk0wZEYsIpSWMNMkhVVMnjvdkLw+ecimmrRYc4odgAKL1YL5/9gGyEoNbtyxU++FNuvO6VZ2B
0vsouxw2J9IGE+2oYOagnlRlydPfgrHAw3mrNtHlgOnl5jO8MPVc+dq9bDnE0I4Gov5vYEwf/IMR
oAp6UIALUEnx0CEES9cG0aPPKkNT7uf32PRp1V7w1adbXb/MXFt81JUWaGA2l0PRQ+5wZwEpjcFY
L4GAGC7VZRoehFNcL8zB9zO9qSk4HtpUmihk0l3M+6AKt4JBESux7zOxBAK8gB228PKKvE/J6YnV
8qRzVFgXCEEhdtvMK0bmYDvfMCV23qZqivc41rtCdt5M7+WrqS/8XMTtrSWZ6XZHv2BPc/3O9yK8
XI2tAOK/abGZr3sDTXSNAg786rOMoggxVO8/dm80dnR0IpxSuzUSJgubpvH+n91gLwZ22Qxbn9no
AmPoyIZ3JIrozMeNGtfWayCrP12uUBsfzkOLd2/DX4ZqBUZJEIi8jMoOyNVuyw5JNaaTz64S1YfO
YjTP+ommzkU+mnXiOiEqEWfT33gNgu9RubxRn8qYNkXmprxKH4xXIcK3tL9KPz+aN5TvW/Uv53AI
hXed+08ms5UmtbM8YXspulgGWpPtolWadHMOjR5YAb7odeSPasrW6lk9wkq1/BgVfBJ2idInzEio
L5QyjA8PXpU0nLqLB/K1g3ox5Zl4w0C2dNIdeOZyHNnMG2yDBwStWoVb3hiIN+hWpx7WvJJ9jIIy
r/7/Uxv57frpPzCP86zrpPVqhjBq+p4XuLr9IeYoYtGyGhNzdgGh0/zZ5kvYNUP+LtCUF7kOApw1
3NnTeSsDNxtExYbhjHYNKLEaPG8Ishfq29gi3Smakc16FJYqfo0yg0X8DQ9v7J3F03BKCXnUKTo7
co3Ad57w15pHvNnieVE00I1GIObt6PruuBVWRtqemq9T9vdsEl1Xi/qTIyn2PgwoLgv6OPym9BGw
I5VjBBUyXR1MFSfh6oNHr6nYroKu0ByaPYmw+LDgzjShRRjpGqRBTY1LZlMbUcxNMDZyVdWCfpkq
FUor4cD06kzLfbZGo4FRjh1ZdItKj3fXd4S/eVnJu9yHbx3KsuomDr6j3P+tt+g+04S9/a1R/88z
/9ClPFoyoa2Mr/YvHZlF4xr3pXYwLtLuZAMODeXgKHRAFExcSWgTwkKhLTISRjAptvGcEjKhIHhg
pLj2ED9IduMNH/278jhJF4mcIjqBNge2Q3TdE/CYsH34D7bX2AyyynazrX4tSQgCXfbGWVAdRm/o
c8/pqHXvABAZn32sOP2wJbKwyYoCcSM1N1s1Ore6h3Jzprd1dWxuj+NA+rNL/aZ5ZwMe+FnCqMfG
H18kW2VEUsJrofOPpHDz3dIvRKvcDMku3L00x2NKw/MhMpLt2JN6EyJw9KLFQ2cbTTpx3zqoI2uo
zmVAmt8lDH73DFki4NmgNP+6R3r6P/jBWdhJda49nU69ZHS1PwKepec5w+hs8jdF4ScKSNING1FH
y7VudXZGHNOmQltAiTV2GeN08a1DlWw8DAZ8zAnKYBF/3Fpyd1248cLPc41C+gxAAGaiqXOEU+1M
esfYLkEEIXq3kreDlmgjyzSlDCQvOi7DztEfMUSvLP6YiMNSsy2CiM6+THq4Fs3GpBsuRVs5WU9Y
WAfZYgMRKCaLYMSiEHciwfm9LLcjLIxrqJOaGmhR3l1DXl/MPwI5PqZUr/v1w5kcymqdZzV91hOq
ytBNNNhW0aRJ1vWQMFq8F1BEYKNSfmkwapsft4PN7lKt/AMQoDsWOgtRrH28MzHMufS++zC8ZEHb
nDMsD0oo2Uap2z8MNXNFVSEkkSrxnb27QRdyY9gvqJ7BENVif7HM3S0ZsPnTsPPtdB3eyKw0unbo
lp4yQOwFzunIghvzJD9nQCGDedERCWfzimqI3YnccDjdNrBzw9aqOyxJrrX7dC5xsgh9bJ5bJTq0
2qNmDkWsAagtJIcJav6GriVEb+HHYR8ftanXmzotEtO4n5Tw8f4XIdG52qyiDwJxVsSZQcv+xG4S
DufZX+T41TfPZ3GAqvLPO8JZqHNI8R2pYjPVMunKrUaWFDMh2FD3SCAwWexF3bxb37+wR5aM7lhW
jmcamDCokx/gXCfU4BwEP5tTvrwfAfAf2Pi8NKtmaIXq5Ak8zAY8/aVEKWOtPlThfIOWDQPuNwMX
HmUoEvAc1a8HA65x9fQzRMI/dL73JIwu2TccUmFHOTyUbJxzoXFhhO4EuhST5X7t6uewcsN9ZqQt
zqWL098u/ySWESIl75Ds/2dhRpTQ5po+oqBvlGDeF4jFfusngiz3vmB5rlpSO4pQbu020ZvGYW3t
bDtKLgH6K7dDLzvAdKGEn0gaWo1tvq6yDJm9W5z+fCNVV8o2//R3/oORZcnkKbkX9t4U+xvCW1Qk
ybItO/0EeeslSrXEipNa2s/QJEGgtmDYodx/OwZWP436PFhIwFANl5RLd4b9EfIBzf3gUBqmqnsG
hfeOb5bymWatrKO5VKQ0580QB6Oa6f8TdtE0n7Bab0gho847FL2nTZ2R39Fa5qZDHlr9iz+CXBoG
LLkNnddBaM62hV0YzaO0lB/+arCn/Qe0sHrJT8OVVz51EZOLzY7Y2xykTFo42Obpf/mMYBKv3vdR
Bi8f6TPCEyIyjXxqYZ/HJsCnSkOPKbYNtF188RR0Xs0QcVVrmr8RMQDS31eAHInsTxZIs6J6/jCm
Ziaj7U7ZJSTszrFNlyyWUFCFumNRg/4SZJeJLZmuGVKJ74qUPki0g0SBEprwhhLFUdEBPFZS6awI
0YKwH7+QJvIeZYzjir9+OszE0hqAhxwgn8FcfAlIjLDcw/FsnsAqWw3A+jdyDItc7o+NbeseDkBN
2YD0l9QqBNsbh7PPpj8Wv3ywlAZBlPj4SIj/eAYoKqgKVahpJCm0UFgqfdtkW/MBUFnaB681Af+4
H87svNQeCFAzgIQMeXuD8YKMgHILo69T2f7doUN6AafYyEv/4Vt3dqMCIZakfvBB2ps/O1mKu+jB
txLsnIsFrBVE+vZOPVGcpvPJjepDPwXWTRLBx0xjjF+DpVeMlL7wOw4KkMSzj2n+6WNK4V4/Db/H
zF9VsLuNChinoUPpxodF3tk7LvIepFZAGzcYVhq6URLUgx8OG6/TtzeoLnSbFdCeS5yS67wHeWlL
MSbH0vkTB3mMiuyFgNnhx0Hxb6c5UJKlo8Nc+MyUatavLN+OBe7VyzcU4jURTz8th20ee/1c/AQz
ylqxWnZCEoQMGtmx/6I8qVTAlyZgy0ogBxXWtfz9djfocEU9hVgmxpc2bfhq8+pc+IN1Rhv2pcDN
8E+gauHgwVLMYXR81xHq2kT4I5iHO+1aIoZCx+kPkcyUxVNV26wWvqvWZTQsGmgZF/pCublel4O0
6ZVsGhOmhxlsV7pXxG1Wmy45fSXqGmoBp+iZBnLsfl/rEna5w8rg16X9c2Wv+Cp2Wsy4+CngjBH3
ngi5UgLCw6fv0QFdl9b54R3rKCaW72N44HyLwShjzuUF7AebigOpMoyyDFKs0SiCKmXRg4kAJQ1C
hQlgJPOn03CkpVyNicTaVjCYvf3M2O7RC9dFUlUjpH1NJtndp/TgfvGr6KMxnGdNbf6FYurRWui/
XTByfMolJ6IAMZSLfO/XmmEmdbZu10FACrcNErLSsSKgItIfMt+oM7Mverpj6pIU9pRex2d4XUjv
fIvu/oBe3ulQOyZAy5pBas+lqNL7A+ZoLlxbK39ODS4pwWE2wo3b9q5vHbIoiGSLNcKIPIeeGGi2
fer3N6AJYy+z/h62oYbaS8yCY0RRKgbyCEEECDpBDibc+u9t+YHalZNjTmvqE3komxCnDtH6qGV8
STuEpclrKQOg1ak8GIQ27oQWiRJn9uVHiIrvcVyDEJZzTBtEO3ogn3NDuV+mYNg2mWyAmTNv4FNc
OYM68n0W8+k2DSXkgrJyWP8UjmtVpSglP8XA1Mv0cdHhrI+0e/c1CaSPmpzC8LZleO1paAmnU5NU
bFp0R8HK121EICNgMAGRXJ56JupdWGUp2QdZkSRdO8Xzybh9Aw5lnzu1TwgGMAP03AjNbMg17utr
T5hfnBzodGGe8P7mR6CFHxvvBzyNVqwtEhKVv/vp0wH5KzaH6MVLp/Gn8bKRvq4HP47e037n71oS
A+r3r8iZYklwJctq22On9ueuY4l0icrmqbPZMp1DodfV4FcsnG7UJzsnz7seBFlfqVxCRr1hN5Fy
T8no4uA97TD1CxgjXUJ63sW4vj00FJjL09VPWWF5Y1HhMHW/u/bJgJg06SDO7MgIJXcSY62iH+xi
fPCf7oLdUnZzHHYuQxhHyB/xUWvOEkjEkaqGjTRRuHTbHlWXeEZ3UJnjfDORB6px75LOHfsQ/hFZ
IaV+wIZ+Kbwk9mhhhs9ysk7l5M7qjq8X4L6nYVCvbcHUBKxknQVr1VNKyIdfJZ5HS9NX43G7D5nI
Qbkesnqr+ww3Ldbu8M/wvZw4e3eLsCVkMa0q8edk2cXkpovmlKhJ4kL2ARqNZluMCoc+nxDuTYzk
Itcc+Qt8QkPMT/eAxLff/FJt68cXZAMgCb7DIPWqXg8JK7bD9qc7Mizz3R2C8nOn50ZNB/zjtpq5
Zm46J0o9FjvSiD9RMK9iwYrg+5mux+KZy8KFx4IW8GSgl0ZN8wtj1iDbau7rSk1+qW2eEkJopS2t
8W23m58MVu61qfwqyaLxv6SL0qEx/579nUVxE6oWIOdO6o/0UDQCPFHp8CwQKU8peOtEgZS8UZ3L
8boBGV6WkpmNdo6Ehh6s9F4YA1vPW80+1Icr2r3F1SIy0nQR/I3+i5yVilV5Kg47TCNkuWnQIaLG
xvNhA8v1a8kDSttPU3IL/2C91ArgWxZIVVAnJZRy71HSONoRyebrOTGXp1xFF4T5lHhdXnAEZl15
SI4CDN5KbWGmHH682aGPg9bz8Qnluzqz3HwQaXIcXEi3nxyZ+0gtM1Ymuqi2gZSAePpIJpQmRwbN
CcIsaSm5gmqLxVZGwUM4meKytBpj+a5PKP5QTCT7LQp+6qt/VZ1kyMK1xgrhWhUqwgKsxQKx5fns
nFaF9uPbPTSoCmLDqYkJspp3zI95Ji/9lv4YYg+flehalFZPqvy1wW8cm3h463ZZacjycbHGVYwc
2t4gocL/dUQ+KgOKr2/OuvP1ijjy2FOaGcjHjYnLYU2NbFzanr7iIFK716YlLZCuIdZqLJpNRR80
PNisi1Fkr20o85jViegvkBrG+A5mQ+EWIWloTLg9ON2bqAfNL8OIZisD13GN76iCZjovkK/L5shN
1AJ/xSZMyOPK4S0sM0HFHBUG7mIhG2ljjmJP7gV/pDKzRk8xjGMy1v6orhZGDoB+8IO0jQKI4Xxm
5qOzsGuvTww6GV6LSf2MUAjXgto2/6svajq7bkrj/4gXyLe0+x5Ova8nBVvTbIbTp6lI4LL40/yz
PFNKZqWU6bbB23zDGX5crYN0Wj7fNZM4QqFgggnvVt1iRtAqhC1ezLXB2Cwxpz7CDSpPXWSNNyFj
YqpL3Iv3IPB3cSENPvUIpJqjzosK3AR4BHr1jE1wNegU+Bv6sA/z9B/F4Bko66XJKyS4WxdMQC/U
5n/fJK/Uv9EIvaAiWchXKs7jBq/9VIejLxz8MpEiHWGUqTkjtzYepjmF61dttHoL+W+29yVCJ5hs
IPgQIEyV1o3hIfJHh6kSWgLGXL7bAx+W+/BKoyNpgt/cB/D6K6aMkMdhbLR3hWZ+Gew71KR43yXm
0cS2SAraYKw+msFQ3fxneypecSdq/WYoE7GU1njMF6JGykOSs3wiilRbY8jlwL6HFTSx0NH2YlKw
1cPI9HBKsALJ0fbAqSwGWbes26rGm91U9Q2tgdPKTJAM+/bUi9R1nIyMwlZCbqN+l06dnNn2uH1T
zm20kAI875sWu3QUfPuLxpc92VHB7tNMEYFOssqtwAhX7iLcJOSHfeP/FDqBq1YdAXqQtXqDIjPY
14tUOar6JY5TH95tJY2fejtGjx0FxNr7uBSZCHCMK8Y/5uBmA6ZCDrTtqfI9yhxyEwbGuy3eF2F1
8rzgYaXQ46IcXGTrt/V/O2HvBtIL/IEBrhmgCmDnCbADDTcUc7ZEOhQb6SJcxQAIfAfX31+bURGg
YgrLmSw42rVQFBbWEZtrj1K7xhZwTx+lG/bgiC+JI9md9xI2Hgie6xWcVPeGJHe0zvl1egGwkvJZ
ku9oKc2nSryHCP+aV+pqpzw4JZgyoleQTRX3TxMHPpIMcEQK0aaqhJbAnZqSpRrUPC5/v2j6pC9g
WdUwK/9hdlNeYG0s7qb3OSTG6n0gygmOM+B28fv6MGm9Ic24/6DtHa89lIru4ZWUULPtIc+boX2y
JnO541aQ9RJgcEjgeJ/XSlaYobaeDO79NUvVFoTptAubAmqtT10X+6T97qxXkJdfd/lwHwXdNoPS
jAyrhzphZjSh8Zh/vDQZdnDy1aIAIUCyh+yhQnDLy3zB/gYai9Sqz7y2vhMlpuTsFdfDEmKUGZR3
9j0qJEntU2A1of8bMJWrjjovcdqGmYUtwLVGgb7OHV/IgLcwBiGsth9MmLfH/6pkJgdx+/QBvUoK
Tak2B77tynq6p3X+nV5GD9lSgY1Itu3+939KuxDPQMJVRBcINg/x6o28l0pmIzQj+1wObi4FvW4z
E1MR6Z7H4w+h60BT2ztiNtHiLB52ZS7Dm02I0IGiU+3pNVTIL4RcysBJnnpQA8RdYM30oWXcBawB
euvcQAspmPp+AhFLaX4vsCbsBn9zuFW4qNcA5vFAdrvjKjgA3c84eBDFJj4p/x0pZdBSqk60dnSR
z8djm5oHuhHLEtNtIV2p7PIUOSL9gBDn2EED5YMUtYNGquXjEibj1txgH+Gdyk3tgpBacYT2XWPP
kGCmsUEzNPBbF1UwXbA91B5OV99Q0mqmuQ7n4aoDL3lEoav4arP63FhyaNi2mig7fe6ePMb0Z5ey
xquvHjr7jawd1lv14gx0ICCKS41Qw7umt/cDSroArWDg+lI9ejF2e80LbVQTwEkeSDI73iAaGSp3
M+0RO/NDOp+ZKmhEvLboxHoLEYCl3PAM4BQdkbFFG4hHR9MdgqpdfkJ4UIyiehgajZMP0bm20f+Y
QBaFm+zNo5qUBLE/B+9uFOC5LJ3BhgBbigzH/UTh/lLRLfw8hJgYKNdyGoInzt2zY6nCotgs2hV/
fNECrALkL2O0ooixgcmg9HJlFjzt8BcVeZZEXhoVAZ+Bpv0tswX6cZv+uf/poy1mB4b3A9I58Gkt
7tbI2ViE9crnpLcNtYlnyA8copns1oP8KYtc9NVhymdOgcZY/vZbg6pJprJeEtFXSWF3gXgtB0Gn
4RI8rE15HH3kOZx6nyurxGpo1hCRgLvCHBa+99DnPVsNEt+DAcsv+Z/Rc+i0BmHAnPtE2EiZyoAV
pD4aZ8uSfY/I3WkQcIIILPqfGt86N3rSD1NIP0LhTav2WZ5DVryV0fJ0Hpy+GrAfl6AD2dxYVu4n
2bK8Ja8pzHpvTCjHliJhd/pLVYxGnELCAmajcIl44KBKYsnTYoZG3+U+aJFZYoxn/Cn6Dh/p4/As
RZTVkAZcrSxnFGnOt/h2+ZRV+FguaEQc9bswMy2tnXakao2ItjOFiETTY06fKaVc4IUVv9TC6C2f
s2h19uhBgypBKC94rLxopypNfC5+bbGUUBCCQYH5b7AgoNWEO2lGwjoc36Nl0jjR5x6GLIJFMBZi
F3UDRlXOwbTXXuTruhdDmafrY0pjztZnzRRvMXlIhigv2vZniGQKvQycI6txa6j7JCcuANN7jU3r
/2Hy8IQPuh3doSEMxcEIPI9qKqDIER2eMcpLVP23njbPREaRxBNVoyOcucNWSEWMqs4mV9rYyxhS
+3VTF6NDctl2IR0SdzlCVf+7mRV+FwKDhsHQe0fcKOrXjip8zt3f1ujDkSwefRnqTLezIRLdO0pc
TaMULVuPUBfWWPFyXdaajxW965HH9RRnmHBpLGDshSYebyQm5ZPYA7TmhtTPX1eKWtgoKYaTRJxJ
Qa9isYqX30cHPMHxkBTOPmY/8yNkE+ajCCtbeLzRZsKJscASB+T8jX7bPvtYbM2qoSjUL711wWIl
8ebRKlKyzTl9wPXDMUg2XYV9HLlmH7n6ll0fuWgU9LVyoAqzOHO/z1otpjU4rM9i1LqTtygZaL78
h7/iN3tvLxu7k6hc729oUicDfbj7aYnQC9qu3B838N2MIXBFNO0hFKDmlobaGYVrk821R4iTAJ9k
vbXl7+CtBSt0i63MfKtvgMhBXBc+DTZF4k+qRa/tFtg9VX1/cRLLl6oUdt2hS8Mtx+dO4WJupeO/
TunYsz4LNHk+qQFmtGMfmINaPAp5xueuvvlxPqWEypfrExa9poYsZ35AZTc6HIKuMf8r36Chc7jp
iE2YdkARvf8Y/SvVh3nhaDIc44g42gG4CO4yhPTRBOu/daSPc+nE2VtT6Lzx+Y9SNcxYPUW3oKFA
8p1/5CLu5ci1Owb3cN1owKtQYDyrJp9OGNq7H3jnmOSyjhIcOW8yksKzgNLlwVGMrki5zjsGHZLb
OuGDlNBLovBjRTtuomJmOxeSfNn2we3KHWVn7SYesViomh3M4dXhoV8eRi8goFYxNhZfTf4R8xQy
ThWGSzxU3JfeQIzgdi3lZNQbRHuUme+VcMQtQ3nZJED0gHr3g2e2NmhBsgsH8hrI58HIU5i9T9ZI
YbTnpS4Sn0izA7ZZGR53NIqccQrdtojkgGeFx38FSN5bwHmuwzhCEQbOimKcMqQrGP9TAWGTZQ6n
9+FRhvmXpz+3F5FhqsgmyxzRgMrLZH/ZcyI/plxmAiHPz3h1S0NuSKsLM3EcTzSnkhlqQJEFCUwz
JMbbMV3I/gKU8KyoavvZ4cv/IhgL1vdxwAMHRwMHukklQVUzza4hZvx0Pl6+Y1o90rLDFXZIjXYt
wOSKbBR226rcA8RqCTHNiBxp/KHxkj37xpxw9fPAMBdmyEvTOwGr3fvdBcFAx/nTiYMcUiGLp7Z3
Rr/fssr19zeUY7dN5oSvuYZaA4LS7grAb8Kpjyp6okTe9MWXv52gMKIA/i5WV3jGvdp9bvkg8y5o
wPtdYHv5LJV9MfXL0RStx8Qqw1f4Cfrb+wZ7VGwYsyQPr2nzQ3qBEuAa2Sgh8pfhcbXu43yzrIHK
5tlJ33jp4njRkbLEjAHvL33DC+R8lTcWsF6/xZFZhBKXbCHPmrSx7Xg5eG3omJiqZ2HXmDwts4yz
xJD0UCuv1p1/KFHT4Et26ABa0kbBHM+hItboR4N/IUtMUkioIit+Kltfcj307JtBMcxkmq9HSZIh
YxWfezd2Qns/bDvf649+uJc6JP6tXE0ErpboH5fCJL7BUA8iGIXcDIkQvtAUwHcPbvlt0m6SW25a
hPWbp+b8YHN3ELQmDKlIX1ZJqGsG+YqQ3Y7J7Kv64aPG0Wjutl0bUO6A6TU9ItU6qTH+/GkFHcq/
q1gsbAsdBe/mxcLwPHUdFV7D+2mWgJTSyZSo/ij1lMCBYbH23rxBfQvwHf2HFfSEN2zmUo5+M8j+
8MQ9dnk8jJ0psOzQoceZGm2VW+ZbLe+HlClUVjzlzGPAuBXv/KZUZTZEHSJql3v/48drP7LIj39Y
2NDsXgrS5mnT57UIlcxk0xfSVsKUzAS7XtrfdazQkgXJ03TvjToXmwkzNSVxHUx+71AfO4SBwNzg
Y25NbSIsU07mjus6YxPSqOlnhKGiRFFPRrAUgQJ/+BL1DnhgGByLPN9zCXV2+qkeU72IbcxnAV5l
Ym950XCYwJcm5GwsP57PCM15QkPoMZiQuC/zHMWIrZHHu/ek+yXwXHC2ZfT6GWUH0WEh530IkTIU
rH9uYeY6F7ldvmdEemyBSOx8tWHtD/18ANFi6WZZEa8jXVmLUUWuxe2sDLManrpEv8WsF3kvaVtW
M4f1kJ1JpYnXyINYMK4Lt37050iHInRMs+et6XT1LCZA0T3QPVokqszFIpzA3BEV7+XoadBoMS9n
jwM8WFVcq9L9+00/qEQxktFbG96glk9/fIKoahtkM5GqXS6QnfCQoz2WzSGvPj24FIj6qqiO0n+t
wEnh9UJYWOcSNWSQEDiJiRxJI9B40LfXuzK3xJYVsuxXClM/0LzxCWQmcAnZjHjtJrCQ6sTBGc7G
uLckVfQNlI6kwyE2veA2gr+HCXPdCv5WYvJJSPHNvWAPJZW9ApO+C1ntonoYHjG81zjduwDHhJPK
zynaUD0c4Nywg21JAD0Kr4h1VFnhR6nPjhGYVBowaFvq8n0chHtjUm2ci8JEJqrqU7b0Yp8fpM8X
HoY7174dUsueWOTY3gfK0fPzryzqWqz72LPcg31R7ixYMd6rQ5lPTlR6VktpEp3WLsD20pOFDDxr
8QFNLVdB+VbN+W8sxpcYVRXx7ErKSze2Ly3+Hugozd2IFs43RU0yXB77ntt0s1Sd3L42KZNm5nJH
xrSuXoSVbI1dq7GYCiYUiJ1c1cOl6TRldAbkZTm4v7yl9Ukmhr7GxNiJRX7kmkZLeV9i05V58Rqw
woiEB15l65sPIDYMl6zq1SVAvEsC1J3rUFQncGueJv/JrhvVmWYCVXjL97Bb0PQ58JOUsfHTcmAg
xjk+DTbYlLnUi1Z0CZQIy9aeh/VnVS8xwGsMRvqyx4DFVlkuNZ1CkPmMqrGTmY98sPvheNybHkiL
FzKnaLNJtlxDrWpo3JYRGuClmKtj170a4yydaJmPu7DI+EnMqi1Qk24xH3NLZvCfhGoy2n/3KycL
s6b69U+Hmysu5kCOif5pCbxwTpIva7010Eoask2LlXqdpa2w2aSmUP5pq/M7/pmBnNeKNhgcV8Sj
0yI2gJ4U1ZILtBunhSEdxqVDF+xRp8WJhPPAmK7FZ/Wjv+JETDYWcVvXIvjDtJU7wtEQe7zybNU2
Jy1ytHYEYGB322EUHMDMF8H311gEu/dbHJOIveA45XK0Ddw8ApHQHShouEMMPeFm1MgD+tUFsEAC
8yIcBUq7IGtrjkY5MARFGsw7kzuB7nWGTSvF4qNORTMfFndXDbwGcf8Og9c5HRf6JU4gzmuV7SxN
thWikhR5AKOmtC8r0aT20CYnrxjsH4MhGX6neH4TiO8J0gN5+m/3kZUIJQBvW2Y0zQAh2Xx2wcmM
Oq4Q0ttFp6f6gf7+Il2UPrlHLCdlxekcSoHje2dSQMtkQv1HzgDfICHxv0ZCqTRb2Rt/WTqBBjVo
6EKQL8Fi/Um6WVMCTQMZynjZ7X1YnhOHDFJaS5es7W+GTqtY/B6fJPqBT8GHC/nhdOvYMF3nZbpd
xR8qB8YHpaflX2CSsZmP9fb16JimmMteVvoFvD6DhzmRZvSj7jVCemPb5QJylNTIcD8Zb6kkH4oi
tDXSJ9HCSwtdIzaGnxIrHEAQ725TtGtoJdn8bvViFaC56jIONJbR5m14s+NZztUJH+gtH7MiKOYV
QmVsmdv+hMcf2+7UfX/mwdFePCDKmElaS2qZofs0/dJlPsCtJXsl4N8jFruWzsRsi1U0uqvz7+ju
FdNSK7ufbmMmTBTwmWB0sl4EgIHP763gy4NYokN+Z2255U2jbpFQycXOEfga3+UEa5IItA/voYx0
IX/GfiARJ1bcQs5UoBNN9mzBBWEZX65h51NYxOh1H8o/bLZRwx5GWBNxzFce8ubPnG6YeG5vKDNY
z3sdKzAiVlXjJgEjJCPSR1lCx3dQMnLFGV4WPPP7yT/LrC0Zxjsyf9DwwMmWOQLeecZHKe6Rdxpo
HspJiHAj8ksaY83Jl/Fw9KlACmBDiMDuKiQQuKSAFGIK8zlrqAZhD5VYB1MvyryOthpCEx1s1qbI
iAS8qDAGlg0Aboliu+oDuBrlaRgsr0hQHgI2wTr50DupfLqxpdNMZJcLcEevtuHeaXxcSKLmUElb
K8eUGbFrchx5vzpsPrjoxSyFJeClBaIBmxnKYdtlnUwlHUYejbR+nqcMKJz7aj/7PhYeYohGonCV
qMu/CydYoSFdz0DBlsU+idorx0JgBwxmTw/ln6nZ1LCQoqhoRVAAU4g5iZZcpupY6Gk3LzC7WQvO
an9B+DROiT9PcAaDVt6euJ9Hazce+/FJWB/tDxUXWqH7mWzmmd1LlgAGsUrWNR7DQVM8svXxAmrV
J6gMCdDJhwyx/ABX/HV3GN3TdrBBI3bh75InxEgPr6lLNWHW+Ob3582Fr/w59A659ou1O1FElbub
kGfo56K+GP9sM1KF4szQ9oMmSEjcjlEKijobkUS1RPoKURq+Xk/7pvbPXxVPz7R27BIZ3dbULgyF
3hFaGnYKAT8hxj2MDFt0i/nQAeDCfY9lCGI2x08tVgNSDDiJnYHe67nh7s/W3HCvQdy6qq80iktO
P4xpAk4Q16vqOIfxSRvVo16D9HpNcszgy+rcli/HSX8n6VIR89WFDHror5Q/znKK4Vtak0ZdPWvg
HGML4sqccZb9uxjPC0yO8vtuyA0NuSfOJgxuVStYrwAqY+GJAIywMZU6NfEHrvyAXyJfvo3jw90d
H41cpWEXx5JIwhxXNhn3n/CqmJHnHQv5rWtuuyiQSuynKGTvvsQQ7r5lVcXHp+o/nEw7RCMI/fqQ
XmC8+Adl3LuYec2s0cA8ZbnlbZfvipVGFUYbE19WFaK7UuhdTBxbB/Ise8gEOXTT4WJMNLtNWoy0
k7Vkf2TsT3XWHRjjT1lPNUFlhWw4b92uA8GBW/Y73okS/NybpLlAuklQ4AuQXojHdbge1NxtpZab
cyfK3Ql7x8JJwnFlz/t2AC0BUkVoHQK7aQ5QFUhk1e9CmSJkknpCIqcUPUjFJqxQXuao8z2zkgS1
dJ4zozewit8Ez8CYvUVKlXMcn5eAPrUZqfpqY+o2Q7B/RmG3W9MOM8jeC9a485DinSWxkXBuLBGd
3Vi0eZ/hjkikDI+iiyC3y3n58cLZ41rSnE3W7Og9WI2ziUZJDsVHxT4Lq3rqxhDOEAgMAsWVINs5
8qVHf5vb8DX/Vlo47I7JdFEp2h9GlWk4D9xstvsY3JY4OtstvR9VwrYU7C5sglnTMvOSfh7o0RaP
bp5Vwb4iDbGuWsK4w5/MEtwEFcfvw8lLW96zQxjLCfORKAtOom9GjDrGsZYV8bNwaHOnLPtRyrT/
lQFEwhJOofBbEPO2XlyW2art89kJC7f2OSyJtoP1/oVRF+bhaafjaz9mVAHN1HLmPrgvFErNL/rz
nZCOun6s5MX+jVmjRaJ8pTBNQ7zDEVW2FKd/yq+LJyLf6wlYpY7+1EKLiLAvavCftO3xaHlR02f9
iKgGvsGPQVCqClxkvBJXD7IUzQPbFcSRZlNwP5YR0zQAzM9ZyGDFAR4D/u9HF0RAX5OF8ZRqNvO+
OD6V9bq6sQgXhv7J2TnmH7PESk7R48n2kKulpzFnYx/BbtHEXS9AynZZCu4aScPukdAGL035jgsx
NbyJsDrCv9qeMKzzOLpdB1XsGHai4of7jH8RouEkuC318lTCs2oDWVCJkjLrw2v4Lyi7k7LWp6ae
ix4ExP9O9JQHtmAy4QcLwQ8EKdAtGuA+//R5NuuekDY72a30EIrGLWbqYFpTeZHMHjAePMKITD4R
o2ePZNoqkObxevZwWHCW0TXLidT8j+knj0HLmAtSdevan2JZaqVBoU/ZLXt6jAc+hNXsxaCTiAkq
1/u/1rGGbQQE8M/K20wu8iQezXOnNwyx2WP0pQk0WuVsboinSyA/e7haE/mwf25agwVkUVZuOpbz
a7za580VPxb/As8mV1FFdCIO9sSVTdHaylxCeUM/53ZUQG6cTQUn/H8ZotwEuLOg5aVzTR4oW3AW
nBC/0Hi5Y5WaYjD9+3dZStBbNDuAuTdBhsLYMOO3FBaMJA9vPpN4QO9W3vt7tf8mNKJHKw5Hcb7l
yed2m5a2XmS+4dw2QbZpYlBXFueSvhO68mruejHDNGR6Gz/LiEin/VI37nofMThFlptMrH4nv1uu
F2qg1oompL+O4lxTA2hviAjKFNxNpnmcqqKJcOKWa4qFTzb+U959exGGjh+X1G+X1N+ntHMHj5CY
4Fr1BEtqI8mEaUUkLjCqrXOV8MPLJq/FMRSowjfELfh+ezhebsjUt6lyVMHllJ9x34RIcBEyO4p5
ujRS4Jeg6lrOI3tKHVL4jtgykhpI4823Sq5oZvdDtM5cXNnlwr/FPsfMVTB3rwQ4EvTzXkUx4bW9
kyS2R1gmsY3Ba5PUtQLxDFBuzUir7e6wLr2wmnQzTeTzGSxEJQ8brDxLV6NLf5p1xweCbIbI5iDl
iaofzbKprTvCJbS9CPS3gKusjbNpiQP3dCBV+VnfX2hc8pHWGuzn43IdXzujabWQpRoxyAcnnUWD
u0vK58JfwR/cr9mFAfYYJlEMobeUowj3q+4S67AKygUV/glW/fqALkqvS+GfMkpnNZ4Nr68k9OD8
XFTDYsp31pEH3d/OwT0qn5vnF5XjPN8ySV2/OISbn/87AvSzactnIDUsDsZp8eZmHYkRkbiYdg9u
L6sILcN7vh+hBu4x+S1e7TxhZYoinK5OemQGTtQeF9LZz7MwYpon61aQN189wvxGI4HdRxP6i4QW
pA67dHojGa9S7U7IaPTpMIHOt2coaZEenPwN+jVjH2VKWtCjsoV2ubyhPZ68z5rHXv3nm0cs5diO
yccE783KUoFUAp3xZAC2v80Oe578AeWV22L9GWoFAOvvbthPg1gnYLCQkiOBm2HIOR+DPhER+kPZ
7lftDTjVjhEkkXkw0EofqS+6EOoucP98AyCjOmM9Px7Ey/8/YqHnZwQPQu5U4Eeazjr6H7lD0PYc
WZK8Btxx0I6kG6GNXuhzn9TkKqqUfbWVylsduiYaEbBhllZ/rNdwlbcAy8JNGO8yKTJuqtSKxwgX
sqXDJI+gFKbyKyTTbT2EABMMip1hbRAKFmJWnCuIEeAfoRdLXAVRQx9x34cbA+1+mN6aqCNqZGvt
iYGVT9PcYTqH3pdWlBc8AYfnrMFdj/IEBKsIC/g8B51TRHCmGG0Qd4GmmMUOkjHzPkoLlzloEjGb
gEi7zv7VRboTt/XIHE4w+zBG3rPxN/+gxm2NEd42KmdY6sma6dLYiGGqc+PkmdU72srYQ/5T8aOl
3XuiBNESYBozYb4vpBoRASFcUBCfY+IvDrND/bA/e3caQS06FQfWC41k3U6b+CHz9J67HNAAWJmP
pGh7Ah2xUQZ9loxE+L9ASK3e/swVLQlm1z6UcnSRzQQvw8UK8HGRrXozvpov8kfPOYIQVtEqHaQE
3arobFWhdcyGOtdVStvzW7JBkudXd3iD+zsex5ysWcaaNJ73hfX7mFURIMg8hZhs14sMCH9yofpu
XdkfHm0jblln8zzN2jvLWFygFy2vKcSReMnG5/uXknQUCxayd4g7Jn7Rx4Mkjiy0p1C6EGp7cDXK
IbvDg740Yhs0wXFXUjWhSvJjW+avCdqpMZHBvpizcac6gBIdhCQqLGzd4WG8VjbBP2oPNqZC3gMo
ppwpfS2FSmVAdWfXwGcra9mZoUQvy4GCchHAVXZOo6tBJkc9TCuWLNLTkcHxd/5tdLIfH0VGBzqT
TfiFcJ47U1EGJ/GcA6kxpQ7aKJ7s1NO7sDA/d4OOWzGjAdfNLYXGWdhunS/3901eCyA0w/EEDugs
w7scErUspU607eNLBPgEY7XO9jp50xbGqyRdk4GuMsKqF8Iu2duc2Nrmi3pPAthXIWNJnbRLhyIL
LHiT0QvaipZ4nome454KXyLUjyLZaGdk7H5W8EFxG+KLyUsi1siukLlWdcdfObA2/Sh/B0Z66Mw6
fJvbhhAhH/fedlJCBQBrRAjcGpYvu9AxL5OnWUqHRJkgMAjGPcCQPeys2x8HtbZa4utEAw8wne/f
sWRuw3DqNycqNIe1+rhlOw9+thnV7AhzZlRU+GEbNEo/ltSq7ApBc+balaajwz8pYmnq3i4D9Y5u
BSe7pnZ7/AhBwotmHXOpwl5eVBdZv4EY1Uxjz8fcIbY/MTsOiITgfuBLJoF9wXG1Eu6bOMl8dPCH
mU4CtB0bgHT3t4au9KBhtrK/hoCCCEyMCOjCC/Oe/wKnyDqaSZE1Kyc+pWssbs3bcqqP7Q/sVpKr
ixK1x99xbIPuFHCz2OFAt0aUtzk3DHaHQRz4Fga7+5gLCdb4i73Ule+42qt1hS9+FslsrzoCHEy5
4TYOZhalqvpUcrLZA2e2nhDrB0QCSq8+2ZQTHAUc1dEcdInrCnKmIsLx49j8B7doxR0HSAi1GDCq
ZcyQAf9IvXyi84Hprzr6BbBsjKecJ1foWsUrqGjnNKpT9Z86w7HDc6BfOEkKJQJBQPMnzlieT5k3
7XmGH8LI9x2FT/QOxSpiAn/q+7nWJW4nlyGjfGW+oAmhLgrkGGZmSfVAZi5riElSTevMZuBm2i9m
o6wjkRdK+3bL2jfmdiR2fGDbzc2cxF+lMT0cVWx5jNS1MBpk5EVLfBcNka3ulabrhC76l6Xq8Stm
dPw8LWjpcZCFXihoxe2E177oP5tsFvVJijVaZ10ExxzdF2Hj1OOuAOsBNv/Kv/xp0Qdds//1R/Z/
jH/rHgo2FHidtrlTg/5/oJVh8RxC6knYlHb6ggcLmCq84pdnipVObkO5sCrs10mDNSEYkQkK0Iio
PaOOBHuDjNZwXd617mPkUWY4Iz91HvpFdbi/J9U59g149Eo1MIGlgAzEme3mnvpowCHpyy0smeoW
Ta6q0hgYbyMULCqIesiAXEPF0eCkDw9DHXYy90ujrIMIPitUgQ5hQqx+Gbu95lyWh7sGIzDvRJEA
O+lE26qRdOA0+xi1F1qis4mtJ7y1dwv6K2wJnt/Qc/cRiuM3Tapt4SuhFCicxmdxE91CrRLrgPJ6
+qLGBjlQ57srYAVMBeKZmxbvjVS3Ji29so92Jqp+K1DJeD9IrwxnHYNImly4qjQpQ80AizitlzDW
A/ghjYHOgD9jsJRoTVIL5oZAEcM2ZyiA405gh1Xq+LQ/YLBJbhb6pDRAipxFFvWGjl5iu2nXFKKS
AOizoXTUsn7zUUUfhYh2RHVpi75SjXcB+16BdsVObdklqalXgNyl/uH+JQOq6FOJao24zHnJYxdU
nH7lnUK/ux/1hftSZw5YQrOim86LDRc1pj8fPg//VdiWJ3zq7i8WW9NVb2cYLz9oLo+itghBuWhX
/uBS7gCbpMs6JkzKJbCdVSWbR4Q4oV1bV/xXxBbZ76ipMk7COLOj9zvCV8t9YcUzoxHge71z3jwK
SjIorT9FAkrT0whsPFRyyiQtqiWSJOoeeR0YHIgZOK7rmjw8dFdBurPbZrjubtlBhXvue5c5rztM
WMerheBrzgSFarcrcOQywpl6M3yJQbctkrnRS3l4qsUS7NHvBGbTj1EiwUcnoxsCZtU/x0Z1ChHj
YqsGziNuUGDZ6DM2c1ZnUuvfTb65daA0jx6/i3DDHmC9J77mPGf3CKpCJWC334w2UNAs6i9G4rEm
uBPmiBhn5VnI7DVn60u1OFmmVenqXwSYf+dFUpZ5oQrnyzwGpcmqO9la8viNW7AepYatO+YKcxSf
i/SmvSyVs/FWrXyW8MRJiw8pzeYeqYQ5n30EGhTonJm5NkVQ5WggOeUeoQen+bhSINPRSQmYr6Nt
yKZJz8MTKMJHwFjvcJwLRcBxNmjwsO+3kH4OvmwGi8UHDS3AyYYP6voSRmAZzmRzpalWZu0f+FAb
394ex9oAbk0LGxldiamkqsuxB+5rA6x4Xmg7Pvu0zXUwNQQF1tvxwdCQydVSvxrHyVhDou4wGdHT
P39nJkhOk7caISOkJzlRwSkJssA8krR1VxmC/47CKBRhYMvfAwwzk7eJ07lcrnOsPe21D+dMLK+Q
o5nsNxQsDHPVgZS09skMAoh1zCaMwKQ//3Vb7QcfWL81IQpR4lzHhzeWATyOxftKzuw/LfiTsIHo
sadeD5iAsC7MX6xeoC1sUPkujLxhSH1JRgFcNN+o3TN4TTT9O+5icTFM4SQL4+sLdrzZCMY5RHzX
wxnUYquqaOAyiH3bc7oGT5coBIhy8ePEPtN0++yVARKmpXfULliaJHSsuwTH56pUWHVPBgINTrxU
Qk0f6U2QxfO0wjDO2bOq9ENBoMLDnZ901NDYd+hrgxWffm+U6D/C3IsrGsfM+tn08hrK+yRruigd
AlUvM7PI5s8oM3kyzMq73TlTDU6zn9AvJKJZ/knALuhHazTn90raOyrqLllJfYZqSxRzL9Lu8onv
GFui5CaiTLLGPMPBgRMLlT3XmxIw4ojuCnGLabEFsvT+d5vBTfAA8fXK7VXhdSPwKSZCs0+d1ofG
Ju0ofMdVoN3imO5UgDF5JAvZCcAB23cZfm8smGzQ/Pz4/qI9zwswpkuk9ZNT9qh/A6Y1NpLmVvAA
gVWEgv744AHP5OQr0+RuP4H+t/ZQSh0fZkqwk8dL93Q/P1pwka6+fb0xvWeyexEB7XtkI/sXymQf
8Ro5XumnL3pSrHNwR4x6cSIFOxXhk5GSNAJ4w5ENh6NOyF2eqEomCMb7j/wgcIguHrrpZ1XPWTxG
hGHUtcB+VsXrmzvMiTQG7j5y/CUpPEyDvqxjdErRItv2CbGbmnH8H6oi3AFY6KZGWOyCRC7MsEK2
YfbvKTxqCYJr4TKOfVK8WtpmdLk2Vwnn/eQhp14dsm8HID1iRuR5YhSPsbaLpxsHBTXoaJPJl7pq
HO6azlF2cqLCyStkU+g/UbwFraMRHxOc9iB3ukGbupQF+i0m6VFeTIb4+vZpa3c62SEU58aT77w+
m+4JFd8mwmoul3QBFe9VC8qxZ19zJXq1XnMiKJquayCucmYmPcrXjq1rf2F0CNS0F8J2nwXE4UjX
T5HSFD3+K/eQFTiAugOVWm63mr5xAlNrb/dHPXf8ezH+orPeNRFT4LdUwNplPIxZBiLHElkL6poD
s5ufI7mXtT8IWymC8C5nh0H9KJezHclUNS3evqJECnH8qbr/Q9rE/M6Q0DXbH8c+Wvk4+7iLfTvP
BYRTYzKqT17N91/pue4QUy39Tc/TaCwgaAVwBkG4gxC5tvDiugE2dOLEVF5ooyEPu41QWCEoQ7Bx
5hbkjxoFIBWeG+OFBsc9YCFSaWPkyU++hgjoeGRwPl850e2YXwn+gZy8A6MBqAdqrOr04D1ImZLY
fFQibA+U+IeuAIQ5B6gSfjvDCej+E4KlyM2yc+5MEiCJ/Vygz9MigMrRUS9Dm5cqZzExOja5iFqu
ymjl0dgv3fATOC7Qu6/ccR1i3g0EHMUizHAJxCDJcyNptM3ki/QzCOAq8YFoniEuEHKOvT9qEI+w
eXf8OZ86NrTEAz6PT6KNfcTBUAUBRd0ml0mk2zf8f77guhf9Jv04VTteWNXBkCle291nzgrXfYWX
id0gX4kiqufxqwZfmeWY2QJnqqZtqY65woiG8R9Cz03yJSxDiW2+CL6Xzq6ZVTnyLJNuqFiGKZgX
Od0NwGi1+3n9hVWhlRK1oYlKBOEjJlFZSY+rZFKWMbxCwv+zzgvWn31nr/usdg4wwmGqK13oE2IU
xwQ72UI8+oaJO1PTirSPSLpa6x5bwmR10e4dgiZpxG6abqKhydjWJUfwxcdzOfRT5iJ068CxbPKy
Nu3ltfVYSFuT+SvYjjv7NT630DguMV7VGRDWKKN0uk3nYd47nC651FkVtoejsDPBApynZc87cczO
VzFodT8L8Jn323uWXbePh8qW2x4xuAOfYZMD02i3vwKlrjuU4Sxl2f4rKTq3L56LV6Qga563e7D+
6/o9ylH+qw8rtp5RR8dfUofvXS574YEKxvcnmVgsZBIsiRZvE/JCsWahmb/Ga94ZuEorrcI/xAxu
O76ZiIwHuc4sxJLsfRQtNTjPWOpdmeVcg6TaKW5DVoz/xJOhwHiJRuCR3XD0nW0JC+MIpKX8QFHr
pmbmmHMHpnMgnYTuk0lUGZGXxxgl64w/cR5Yo6zYO5P94ZGwtP2SotiVdBImg9rMl9XKGlIt4o6L
LXpBJfD8z9h8xqk7+Jr8FW+4f+QM6ZMcdQDRBxtGipqTbqAB7S/m+HkDix6NTxj5C2v6lYULeE2M
1cFelecbp6NOTu8MPndtSSqjACLEfOk0S/d1tkshHRbwumBq/HZjG96UUzpZoR6h7iOUGhDiDOuv
RTUoNEVi/+bdAHE8CXxmf+GBmafzmEG3aMzydOwdUIsW9KCWfuSO+jEEfH42pWJX4mjh6iwTxK5R
Qp0HQPLf2bY8QcAdI8rCw9SLy1Bx3LDlj0zWA58uQYWTm1QxWrEsRiH/tGDHkkB2zlNXxE7Heo73
jvjwMfo70/9mMzMB4lzhberDYCoMaF7+8eRwVeICahH3JhZkT4NesPmPhH6RRrlR3muNBozvz6Hk
xDE5Qk5NcrPL06lLuX5Dv71tM/bGVVbBwnmOE0Lszcj13RyuGnDz2jjChxWf7cPO7mP9Xi3UovgS
jIp3pioHl/wMNZ25VqafZKRs4aAxNuCHto5afnOKpvLUDyPfFrnVhs0OA5qbcE1XcRyP3+gOkHaG
u3oQqgYXUlCwQe78RX2bCbPsCddXTkPDBFvL4VFK2zRkDeYyIYKkc+ptZB3QWdmHJHReafhRUVJu
6bn4IVy77chRVgWwN07ko1p5Yl3H3FPkA6G/JXklvk3HuO1dPHD2pBlrqFbE7zX/jrBw0n1s+YUw
N3b6qUBgXsUWng3k6S+j88pibLcUy3tafWsi7MgLV674gO4tI9VgxryDrqb8deu6feCSvrrM4eFY
DwQ+tnph8nmPpQydNC4BIUS53lYGI1zERu//GCXVOS2BWRkhHT5lVfijGIErW3+JPmGn9hogbOR7
OJ9nNOAnyF28IZt86QNlLe6R1WJvPd+T9AtCW9sQxon/uBf+bcHdwA8soFUXhBGY9RkMLqk4LZp5
7vX073sTu1DX3NHm25ytiDSb3LrLHXesr7/lB599lZBadXn2onvcqOZuXKcM/yUPwezysY9mYY+g
5AFm1mQHLb+t0I0QTg4L7Kmd6uAnb2djDyW+lcw6s3MqGFs11yZrWLRoNg+AadAlxHyHa5nGOPRB
PyM6Fe5ENJiH2ec6z8q6r1RfYu7hnM+XZGJwX2BM52y9Ow1HXV3yL8SNOSNpD0kdC1NlrEN9LqDj
kla3EG2eeusDiSp3VdCtm7WwjxQGIWPLew+0Oz+gyRYpHs+VMNsfC/tM3YW+IogqI9EEdFerUeWP
Rws2rhy3/tWTNZ68+TsLepcBzyw5joSNwevQCJ4MAIW+GwijMX6RZCw6uy56q3X3Y0lwREIv8v+Z
+b1JfYJi85nXSZXqwi0eQXlmUWEXIf5HXpR12uHfvS1eatO8q8dmUepH7ObFgEfyqJkxxQXTrefy
PhTIrxLP3n04Ev7kxNKUNnqWGPZG8s6kF32tdnlbslaXdHMwwVJ6/sM1I/HTPjYYIICSwKIKsk/Q
ZxZNxXP+HbeTRASgPgs6dqA9oe/eHwIB+CP6hFadVWUebISeF0kEm2qjkJiqWUuoEJk9w8YmDTxN
fyLjymC2jUzXYvPdmQOxu9cRCsdarCjHctwz/YBDuDy+aCSJ1iz2LcQlRD4ujiH6crc4+0UeRRxp
c1Gt6U1od4QzDTiE2dUzwKjj/qaq4Ork+cLbtqXky4wXXWEwsiI9Z1ZOm61t7QdUCDLgxdXW6QJe
q70bNfUxuv/+vH+3azMb2O0sWbR/+O1Cs1L9Ck+JlQzEQep4dRcNH/Pc9zs1U18ia2gPtHjV380n
wCuss+HFT8U1WWb78G0MQYw/09NfvpUlaw00+N8j2H7vRFCd9Uvpp9xRlCAloDEeO5KcDmlGWkOI
gmywWYg5PGQi+xu97fA0NKSmgSor4S28tJRRtqWi7GR5niocGqkj1+PEnoKoWF+kPMj8FHSVghXW
CzUYECVo1kn1XTZPu1H9nJLjcDvCQgQerJ/U00CmwOKmcKqVBeHZCNXn0xE7rW62dTliGkDDNKsy
yl+rDN8aIE4+lHxYp2m84BIsNmRSpN+FxHHGd/j7UlQAI2e2pfzKelolRbhlXa/zD6D+l4JjTEuV
uFkYloFl6bbeQ8toXRacReGo9+fTvgCCPOn+2NqGa/oGcDcHUXu2psumctBrlJ+Y8bb5dA0mT+98
lD2SBrU1cPo1Qcb0UZQmCkG9GEjykv7TUbrRQydbbqYqbUldQuLbYIoCWdEIiH3Q+6L0J70N1S/M
MIPDI9dlLdQyVm0qCG9s8vNPH7qiu70BCUhabzM+ShRpuLT2dvuODlReSGT+7fzasN89JxKKfUhv
aoGoe9q9WSdk3Lwg1LP3dX7mN/INYl/RMJAYRzmjWYdRJaXRep4kutcyfdZcBj11dJ8CYX8eFWxN
9sc3/G4GcOKFiUwKpIj9wMHXkBASO7NjDChgGuFdaSELZfC4U+pBWWTV+A5YhaoPbXeeM58a5EHL
ZztZsPVHksu48Z6w2+kE2Jmf8oafBuMYu0Jey6FmRPSziPsVOE1jIuhYdCQEEQxinAemdTf8B62d
CgjIDO57kM8QSqejcjJ+6pn+vpj/Y0W3OFcHP+T6ky7nbFWbPC+brjT0EU5WfTOWoagWCvq3KeEO
iN1ZmkR2c/jDe0iZttx5wxi5LuWk2F30xsTXmcs0aBHrcvlQJ/JLgy5ry1qSCEobDRFjb66UBfmn
oN8lXe2tOAIcdNGTPefO5b+0gX35SvvYscBpgu7vi8C7XRmxnXv7eYY9Qt0YCmBaF+a8jwFSljSN
9XtQEU0bNUtIffrI8tO6Mc7kFhky6SO6xgRbWQ7LO9Wj6q9ir0G5hmVBzhaMLUESlBf+s78JFpgn
9RoT9AWqE7pqzLIf7ZyEiALsTAaosUwurTgXC/SL84G7JADQlCiMyxR2o4t88O5VsJgsY7M5PN1B
ksMu2AErJqz8psmPLTc0y1Za/AYuhNKBkB5BL5GZZhbuf4u1q3uChqmc09GGVk0RsLVQCWDwV9R6
tuSRe94zApcJ7uGQA5pxIzfymRpOLd5XT6ZNALy4zLCnV8rN19+ns6NZaHdbiJwpmZKWHEg8AjhS
CS3auGT3np2n0ZNiPYs/eEY7auYefu9aL0FSM2cwvpC+quLBNAlk25J05jj/SHrlDPUqgJpSoj6+
3xawLW+tQIvnIgmKPf2GPxMgZKurdweDzfebM0XHhOZSaUbFfXl5wm7IxCL4Wah+xSB8ucAyWAb6
+RicZ3X86PniCEEgl3EtKCXgY99S7QuY6Ufjmt/FgSYdHUWozDDXHiT/Ob9FVzQrRjqO7Z7RD012
+mLvHaika22uGMyXw05d38CwibV2UnMXDP5Ro1daHIwkvuPNKGLQx7lnsqbXTZN66yabmqwx4FD2
s3vCyYX5w/HYSNI1a6fglrnfZgZMZ/5hPEQ6/Vc6IVIshMJFKyD/VMBNIKATjjpLQISGYpNw7apu
265s8XjPdUNZiENBh42LTleoJrcUwcVp9Lp39uN5CiHFmCjmWfHZoAU3QuaG/bZKo4Ca31jDQvsN
X74q5DX+M1RYNO+TUaLnKNrUAYlGWIZrfuqXGsvHvEKnGBX3Pn3GuJtvIol7wDN6ZAVF2HUtIGTn
wAzA4sSCv/8uIbRAt+aG2MnWWV3eYGk1nXhj93x/WrDx1Tk2sBWthCpEKj8HzWYtXEoRSh3HZODc
kNozzyNmCd/paS563sdMp7sYUoXc6YMJzpjPr42p25SM2uJ8Ab14vTAk378zRpFVQmdw793SzcaS
QlKhFn0V6makBSC1LLAv3Ha0XfXIQhUUSQzLOoG/lEV2J81ZQqO3wJ5eH+hGLVCTb0bhOeIe6JST
TRVZA9vjrQQHtfOsr6033uYZ/wlcr6DTrML0xf0JtkHvXbBc9VSIcK4IqF4FXDeIrMPVRwENX7/2
2byOK9uc3btwYJwsx9SIn5reoCIe2aQk7ajTMH79g9vHbTafDUmtUSs5P4ExB11IHwGdzH7LRvz3
A2m8xzkKy40EiTORkgpNcmAKZio2Q8YjWyMROUuLDaFJQmXq4ldoLnQ+o1z+r3JBG0+9ubuNctBy
KOOV0Y4VZKstPtQOgxEr+ZqegVxGNNmrW93NN6cTUMVyz9IRLVSmwE2We0tgke+oCU4/1tiAHCw8
P1dzb1JV3DDflaji4KsIRyGdfkgEgtvkrshi2jcO2HHBfEoYpK5YfnOTqbjG7OVHfudRtE1j8TdS
iQjB2kWv5kmAudu7F1HDKrBBMy9HMUURwVWqBYtxTdFBu++AZaKpyfnPs2WXIKS1s85qjk3mM7H9
ouS56QxdP0kb3UEhmtEK4eQTLwG74MdplBVdF34k1J34f/abysFT2HUbuHo7kwp5923pZrIJY2zg
FRKRxvAaHsLu1XILOXLTKMmLStN+BZK/GtfyHO3jKfxPnyQyxt6K3C5h/rW5tLc0QE3J8EbihUJN
/0Irvs9Pie1u/cg4VATfeoFdm5+aSCFz7bHPiWvY+C8LEJHykctrqtG5pRez1eQwWyTUX2sJJu3v
Pt2ypvAiQZC5fl7dLOuPRflxNKjtDVblq3oxb+94KPM4UAndGZryCmNwuC0ci2x2XJM8rtRauHr/
Ptv5v8p/0LTOE0fdO20FLGjeJzJl8pGCRwxDekWG/vRC6NKCCjzgpa19PxqcFtZ2R6tLbMgWlG1X
lb2RzL5UGPgFwGxJ8cJeSg1BLyVir42vOOwcn/xviLR3eIjRp2VHCRXAELSinmyOe5f0wqVRzqIa
iq0QfffTMmrKP36tCsmoREF3A3CAA90xvdwLlB2mxyHdBR8FuEdFAdpQi4eUOBacDuu+2msPhurA
SMHeuILekv61fF8pAA+SXmRXKb8KxGdQCEEsDPlEcdmk9Y/rR43Zu0X9ipZ6Aa2USump6MqR8heI
OJjKxyfOwGk2VI7YfW/YBNGSVSEzyVQjl9bPTVcBRzjkcYMtYoncvD460om770lcthOUHxIWFGSZ
GhOFmxPqEl38mUu7ijZBOq9VMnksI2C8/AtPgQAlhVgHpP4rPx2kg14o5QRRGkYb+5lqeQRAlonN
8tS6HgHT9nwxJA6wIaDcQHQVF7CUZ0G7NYCP3FelBd/lfo8L25WO4V95VTm8mIP7lbTDa1mNRuiB
GHqsflSBL3rHvsSKjCH5PSNSQwo6ZuqqF6UcSAdoxu0qN8SM9B7AiZEhRVLr9oX4DATXNwewbZDq
CcT5IG9lYAlGk9OrEYwS248Rbzsu0UcwZWAUwnNSKHWmVSf8awleXlho8ftZJBdqu3bXGa6jk/Oz
emprdII0Ss57865m1WIwWP0uJE9cTbUuFE4ytcKCxV7NrSBaZDsu19YN2VbYQPaZ1eLkcQysDbSs
yO5tfwLDoNDnIaTevOweTsA8LWz8HctyLC8oPbvplFSb3dAjcViAbLhLEhjx548NqSDtWLkjoFrM
Cym4T5ycyv/scJCIXh+KZmVkThCrF2RxhHipaQVsJ5r5RCF3G0tEMCgVqwDBbtsC1Dkp/xxCBiGw
DPagxpkqlAnwfQ0xwCqnQB2ZAKAoT3a4lah4aQ6N5YFEzkMKsDuWux53b/kOY6qg7ksDmfjd5e+X
VJxaHmsFXQrmk+FE9A8Hhfn/6KBehBBolv3V8fj7NbBXdgG6vasiOljZTBauxWJzwkjNANyAvfNo
DqLi3XECxbJYXSk350ps1YL+HNGgBWt4oKlN9d82Wz6Up/JI2BZmCX+nMSp4RpwdNylhhWgxXLW0
kEd2X1O3hf6NkFl2VL2b/rbHe30v0q7YkmIlHgxs5uP6t2E2gALgmbBBrx/Iunqp9fflUteaS7jh
ZOlMol0El60eqO+EdpCKJt5umwcic/5+m5Kufg3lo43teqa4TMjLk/rjp7XeI3gYIInkGsn/AgSk
wgTpuBo5dnOD4GRpVV2xKl+cwlAKqZMEaSI0qlnxigfaeWszW7iHKHbhOcij392ZC7V+GckAk/j2
nqiX2yDkLH/EhPi9m9qd2+SagJH6gKK2LBFcv65/OG3zJxuLdGtLdMPKSX1bHuwhr5Tj/pr6yPl+
OUrqE3EG8rIOGN0OVzRdMae+ucBEzBOkCMM45yvPv+2riibZ89bCagcZ3JiwEHFZTvlAVJFHViks
N/oQnxXvKYL1l5SKxO6SjwVsOCP47ZRXTe7vL9JwjkXb2vqcGXn2R8i8MwLdzrGb1Y372AkKJ/IS
v1p3cR7bWA+0v3+pyDmpXYEzzvlIr91QnuIjPSQeSf94W4l7aDmesJ+iBZBD4Dcq3CieYargeKK/
O+n+I5cPU0Mmgk/i4eC+itnm6qRRRcxledvUsle//WR1wMJ7lnEQ63rYHX/P+3L+DoHki10gyqLu
+wd5CO+GvC0prIp2Z0d57JSgx17aUnkw3D2hC4DTiynF8hwzul2JUd83nAWcq/dVEGAHPhIO9M+r
avFCy++oTVFffvHg+2sfSV3viif1ewmVwcHJ8P4ztKT19xeSmGdesN+inIEB6qu0pGRl7S9jy84L
fzItBw2hk0sIErRIghl55VA+xQLjbMAu7t2XVGNk5npUIHB02zEpjPUiHZK/1ZJ1MD2uQuGdURhW
QD/d+M2uO9qp7MboF2LEYFoKj44mVePnGrQ3YuSmr7C1YbbBBxDKEpDnwavTpVW4cT7EOlUWK0am
tdBDpFiEA9HOCUzyxWesk5vGPU1qGezPIeSx0SsZfbTHsbtmc9R0VhpstkPiM7iglCcnMJC1nxqh
iUXp+pEouMJP2UL2YZv6RTQPUEsq9Lis0OnU0rRqYWBxYitdxXIq8tg2VyFJgf37bSa0Rz455uLZ
nYMFjbpw9BNudXvkw2mrZYpoD0JT4qXM8YkMMgEOvvdlOSwugY3D/nRh6eRDTYW9Aj98z0S3bvAt
y2Y2E1d3iErX11PvgyYAqiUAxb4ZdO0bqSjmsbdAIvTAQ4GkxjLiT7MaMAlSQtKrw/p3C74mKb4A
7Fd0ZSI7gnmticgdLNoXqxgLmrprXMfz5OmdcLYjPKxsK+/K0UhmeFA2xoOMxcI0QbpclwG8cicL
3zJJUtqHYZ4sRRcParZGK5Hh2ZMNVAMlZwnV7GFl7o6CUBzFPpb+bl400olr8L2dp2MMfv6LEE6b
hXzzRCd1NQqyXBSsI3RUMeqD945LIy1wK+ObO+KHbavlr4XoeDewlE3l4HgbTe0JuJJoKx1TtgPt
oLlbt6EMnZOmfqKNpR0tSEg4ywAw8fxLhf/nZPoJjLAEXUx5pZAnDEvEqspd+4ZVTsb58fM63Ydg
MhDteu90dw4/OGfKEZ0miwax9msX4kn79EOrb1D2ysldoxVB7D9g9Mo4oRQDeXenS+ZuDUrB0lY7
gES2r5PF3I65QWzqsHl1EYxtU0ySTy3oFXu8eunJbEhfH0U8ukbBrKKhwWXrCx1xcmHDOvtaIZNS
orGkCx0833vzLh7UtK7SH6cg9BxgjxnpsYQ9DwFzXQLFU4qaEYQ45SGcohCVATs8TLKRrd1fwBHk
BJaQe8Twh5mzOUhYRfvYs09vlKV/k1EPvjRbeKG80nyU4mDl6r6GoZ0/uShPiWA5VTHd/KOaQKvE
eUCcg8BJ0M/RA5t+ZnZL8M1IhTdq2qiCwu7SewPG9yslW9d9ytoQR7m0NKPQrbYy6pCjaKCJ8bJv
R5tqmFoBmZyhh/iv09WfIUC8nqWkJwDve+eCgGptAYSMbknn9DCgB69BP6jcq7G1uXbItWuLPxlr
1mAWTZc2drZCetZxADDJVNoSrpY/s67rnsgd6N/ydhRhDuMbBcxnEYMB19/6qBbtSLBmTVcnziMD
NJZxLGvvv0ZOOwXSy4+N6yeoVQ/l84cDNd1sottuf9W5mRi7TZeMmYZgKZuinOScjNVerpYut4Ds
mjOEExdCE9rNeJ8a3nj40hpJBENYCb4TH2b6HI43aefo6/7sYveMsGeQZ90+vfq/3C9LxDABEWWm
XPpysHfRyGxM/unin+rCWKT75XcDFInvh3tfOyJDHanwS855/CXdZ86Vb3PpGyj9gjXsmT+uI+0y
kO59z/4qcsJ1vAHDTCfYJTW5N3OLvTqSdqrowUq4JqRFA/lLjiYpzLzHDsAXTuTpq0b/ul+snLh/
FvWNsA4CKk//fSVthlF4tezX9MZ+vIQOGOd1md8nzETaPWr+FMkDOJCxqCOf40zfnF7iklCEGjeP
Nrq6JgCCRFhNOkuPqMvHXlYmDW9VcMVLGlrwCCnrUZDFLbXxajgN4v5KwA/RKaZHMK4D88Nerj91
Oge9XVf32CaDT8BkVBVpgxThHVRm2Xvm9vdlAak+PoN45fvUiFZvjyW/7uvi7e4De5lRrlxXn6zv
nHSTPl++shrAKaLtnYVLSzJHxgOfjhWMCKpL8eyCkuOpGH1YEoiPJ2ErL/6MPybnLnZdMWGYmtcP
sHymVE643qzst9pDqzuQHmCbl28DB3vkoOhd1AfW9/IYKzhpyAPQBZPcSn3RLta9jffaAlUrThUY
wcZ1pSh6nzrLUx5GwQMU6q465DuyoURDQYmuJ6xw/32d1ib15zPbxIr5HFQc2yPWZhaoJgBzYRBJ
/RYTLTRGc4vBtopL+m+s+74Tg+4qHwuHFRpa2+23dY3FJbtNt6cA5DMKzwA82XCDIkiVFqOZKUwI
feIDgOENslkiBeJnO3zuJKLCE5JGI4KDACKAH2bsjeaQA4urXvOpasZ6NwemgOzU5Z0DAw3J001A
28FTJ6jh+R34p/blwiCZnY1a3vUAHYfIXGnVomICOBmFM9LgXcBtXopL+ryIkgwAQbC4jadZrwYm
yrQBE55LezOkBECLWu0F91gXj7gKeCAN9xcwa0pEmcUS3weOgh6p6lGMlcJdmfS9dVTTP04+Mlb+
MnYgrF8rASlJlCFBW2IVzmVvONf5YGVFMLED9/JBu79QdMpdLCe+juJH9pxQ5M6NPWVblfjutWaj
zE6TminkG/MdlhABTyVCU596Q7LVX6GdEtR00b/7aQFICH+wL41pdtvAYPRc8eQLHAcDI2NPrtsP
s0aliSiMieAVb7LLEB12L9WppiXn9oNz0zdNfT5y0ZklLBRsK4tewMVoW3dTpy8Zv2jUdp+7jZ59
luhJK/T/31XEDnExCcCXaRRvQJE6bZHq6W+PHnIig9HW7hBZH63Pn3v/BhvF8l/YRILcsVnsh8p8
xcmoQOzxiwsBUnsbnyBmgjZiQzBgxgw8L5zZvqblUIGr6V8cl/bgRnKn5aRf8ksqMEAQHazmypvG
yreZDn9dcshrk9vI0UIeYquIUUN0ci8keX8a2zbj8IHc7axQeoV7t0gM9OXUIjSF6V4Db/o4PweI
jySQUNOJShWx+VKIJrf06RXL190COa/+sZEXXXP0mUUEYguhHMl5jirhojv4nwFhKHjgn8y5Ukqt
gD4DXVPzE0rUI0Td6Rj5EENvzR/6fphJlO8EQPVd4xf73BfLRwjwUuCFPqdy99o+i5xkP5oiqF+X
kiYHCBBGCV3Wmk4HeaS42ydIGUL01RxxwFwbMoSzdAp91s7ESgDrDV9kMQCMbvvLoHD8uzBIh4Cj
SLQq3ICPyM4VPMPL47gLw7V9wolxIk6J2TGo9O07vHpAjBPxfUAdgykz41gTf9wfhRb0DL2jGfJN
waa1Vk/oo+zhPNhrGwTDi+5eNo8QxIo4oIOqrHMwGpvkx/OcADbCHQuJrMV0qrTDFmsxh4NrLpSA
a164ebCIUhAdzGKZ+DxMOTq2GCaKeP0P9hzpI+zvEfWA8rdXAHLD3J6mYTNSsJILeypL455FDoEC
lQRdCJ61YNFmWV/KJZj1HXAsNytFAykBNynPkfkiKyCnCXUeYQN8GdlU8CA+JeIeV0Z5cZHO46NT
d0SuuYeaOUTK4pxFURdaCaSH/4EGzkPugsMqiNuU6oNg1X3IKHPjrRTrxac2DvU0MdCqYfhQzkqd
fOzdjdUqqZGnXkCEgUc9dULXwQULZe+RVutQtQVrScoOETp/QKKGiWB81ZLDZ4JMYxb1ZTqh04BV
onfhVldKeb+LMuyX0ctJWRRNY7OhdD1UmubpN1XgwdGLbRk3nVM5cbNarK3T7qE8vWpq3ydlH2bV
ydLKEGrwpZ32tJ/FRbzSpZJFJeXsZJlfcPcojeIOQuQNpyGTemVCc0CHLelQZ6oCL1lwoIexBaOH
QJLkX6fkb04AVgNtJSeBml1rIzNGlHdOZlU0kQyCjgFIie4E4vLuzI2CiH6z+eFoS6SvMQWr8oYL
QtC/4JCwtPyt+LcpVTTFW7c9BzO8X3C3RHJTUKiOFQqnmU0vdum4ovJix+sYeZTBoIqC2kClOele
VSKShfnRFoUI2uSfG1FRQ9mWruBK2l9fA5gedFStjAlRyD0B5R0hDT+jLmDdZ5kBQkSt08Be86Rm
+FEq+tlmDca59Q0VloNU4Hat1JWIoHFo3CQWdFWWi9ARu2zifnoVvI6quKcMq74thOOVu/wQGywj
x4VBp70niAZ7wuqnvXHeyGA5ozbSvcIEimduihdHoeiBeapuEZNTQiJfiewTFuHlpCs2n5TmyjNp
iBTxB4//Hl+sdeBwj5g7bdTLSxTLZVU/RLIW/hH1HSvIVGGI9qUFSqNABrOZUu5qfXKsJSXKUynI
f7aMXODw8AgSPUjiJ2bcIyBdOx7TFPX98Tf/y7UoDRnJxGli2S8i1Un9SbQwvnppvTgtG260aymN
KclhbeDrNNDKYsfIDaQsCkvjVoCHYdrYpOSYWhcIB9oAig37/mfutRFVB0EOGjSKBuS7mclPeLVw
24idmP99LQrdEuS+273arPM3MohBonkxmf2X3Eu33V0tJycQnH09jYw9r8K2v+ZT375h5Or6io7N
aflMPE6z8iI2I5a5VWVy7g1UYWcn/8cx29OiLH+5WvjK9xJzN+bMsTOlos/8WLotcofk8XV0tR6c
U4VkooEHwgJJLU0oJcPu4C7xnba8RrD/fTqNlnmO9tX4zNi/CLoZIGhzQRQJ3SfQt9aAa8XQInwR
4t3EsXZZgPVP7WP1sQUpce3bQvkEwUxqz/eRP7ztog2eT7xfphWb5vXSULTbJnVwN/SE0sivznqN
IHnsIXuYWGDNHoLZyITrsJKNq8r+5LqThsUTbup7QbhEFEZq++yPvAMCfeM+27zt6zdrpPH0bPk3
Dt3BtrF6+31CJCngQDJOfaiE87WOBPvg0xj2NWeTFRqOniwpUetEq4fCXMclGD+iuCBTX9W+Ch08
Q0VVF3f+E2OIVHsI3EO0M8/ipjoWto9itFhzvTzUo2NqPp+3fMVWqZVJKmlpmMUu5BIdRdjWprkU
P/pEy38yqrBl5xaiIhYN97CDcnRD46AoDduUYkGK/VnbXkNfR55TA+/bXCTtPRj1H6Pa7HMmFKh3
3io5TiQE5/GpBkoiPul0bszx77HNB8VQ3ZYSMNQ3fiWyIGNNpUNT67qDYFdoaJ2CL54BvDzlfwDI
lvSoZ40yxpkAbZkRwJxojI5llBYJdlsbmyxFRRIT7gS5C+9NTUHfbMtlKuTrXKyiaGENn51ykcgt
h1zd0bC+YjJGM57FJJ0V/8pOUbTC4nntK4J5TOP3RywPEJfHInPvyuz4PMrg0PZ6y2em+u17DMUy
fhhIsX+j+/EhwtOzbZT3SWzfZmpkCkYz0oZvkHR3ZFhxyMwCKTifFbAxEBfLdzMx6U9bB28XQJm+
93yrH7LlZELrRuMnXrkxxQWYPFux35PpgYkkqKl5nlvJWje+D5LMGuVdoGvITqYzJQNtygNPSKnM
d6gfS9DsPjptgLjVFNIRg5rt6YKawIWPu/QQ10vbJxwAELovgdhFVWIXmkgO2ANxSm1p/0Z3Mkeh
DtRb9JtbKi5PKLzjfSw60y/1V8GcLWxXJ+ChxDUitBGVV0vTJP/ckGrldftR6KLkoXbtFVFCJ/xe
7cY3/xcgd2jUz42jtLu1Zp5wnXdx3/92X9bHwsD4E+6y1FrbO2NsWy82zsdwXcPxpC7goMY4jLfv
TmLe0NqI0gqtn9e3cvVj5Jje2mb1Z4BT3rMfmQQBv2FU6Ra0YHA9v2USQ8NLRRgjC13gNyVwczWa
72oMTrSTHurq80rcrI+6UMC47JwSt4tMDnoBF3h4/RssEsMUnUPMDyyrByqOxvXL/G3PDBWf3iTn
nmrOH/WNT+4YfS+CpUZNCxA07+tTUq5bXiFGDgL5M4kFuFEKuGLr4YSocwGOcqPt1Kp3pyMyLfMY
+gSifp99sSMQ6DuFBRxElls+KFGqIfmvw5oCj2yNQGgJY2xaYY0czaQ6KnVUdZyZw9gyD9mjibyT
WEh51kABE3il19yUd1nhlK9UKkKIJ3am1kGC6Q2hNjhe/kN+o+tL1/d+zIUdYNetlmU3LqfQA25N
3YvBSSGN6bPVYVV11/5e5uU2dxYaqNb8vAuvcvzkBZDM9b8s0udZNROqaPnO5tGk8lgDgPsARgt/
kMdVF29VYIHm0yB8E5y7/pbUL5ysytW2pit5cVrt/qZGdlm+t6TIULnVKew20kYZCOoFt2/CtgmY
oWSqPKfRT913SmLopo5OoLT9ICqSiBkVvnVYUBuvZEwXtJwdhvYHBzdBN4H4/mFjH+bGmd7x5o7o
SN/LdEVsEXTgNZU8u3D8XWL9Q0cPGdH8BNMtLeOTmhfZVlXb+i9FVTAIdGvrIuinPmJMFzYZUv/w
vLosLwh1VH2t9mLGh+ibL7m8Qm/ONXPzWw30PWuzp2B8XC9HO4/vFFF2cTws8kK5tj0q0erwS+Ec
lbsi5mWqsLnVFJWlxqxGX79Us8iN5Y+adsDCky4ju2QYkHZtr0hwJ48lSRg3IZxRK7bU2Ru/cLBd
TS5R0KEbMlPnOIJV/woC6GXvPv6i7/J4cl7f8hR+ZSTCzdw9i5C6AO5yXbQv/ZapmFwQylZ3ASkQ
NstAryR2VIkoEwpMTARsfYpurzoVECjEg34IVkZINwMZs17fWxyJnmX9nAEaOXk57LU5qPu7tZ55
cqUL/zwElCRiTltZO2EBOH0Qmj7q2rtJAwUX77c1byjU6ZtxrWmsaxVIrJ3kVzGfbNRja+ED0hEq
OYRbaR5ahUfgdNGoR5olrdGO4rakZzPe2HYruEi7EeHQoVeJaorrV1Ie0vbSxnigWNEmmC9qDii1
QRWkVkSH2ql/Uyehlew/YwFdIPWNiB+7bIsgDrYSBsz/cbh7aP/UJ6w7APZtkUTxkWArh8vPCV85
oWkVKxZtFNPfTtJJAlpRLKi/5R93DtbLSER0DdbGSCrvlNmm4V70mvmTtS+iij2mHE0GKELbs3OA
PDcvlKLaYSNijPCNc+XzG5g5Wg7rterPJt6oWGkv6QJ5e5krKddnbuT+kdBCEcRt5UVe7D8X0+Ia
d/6Ucby+LKFV7pIhK1vN7HaER3R9eCXROlMhNudLYMmngc/FU/yJqvOdeqakl+m7t468rCkaS+X6
VUNT996oJ9JGiyjggKp7MGOdM13efg2FqNHKWZBVWyYNY5fgepa1hp9s0Va+8xqYeQXM4+IPc1Pu
06UoqGPWWJhHaVcgn08L7UiRTPEZt+rAxhQUmqsZbBy2d+QeIA8eH+pX/k8i10HKZcS7iAcyzdUO
iNZ4DJRzwyEZNRQyGj99z4WUGlDajfYnGKBisVCvwRFQUqRA7mOX1Of0LYgLFfOB34Aazg0SnBU0
2qBLNXolCxy5YT8paK3X9PGlgTqyO6aeKLfkm7PVgN5Ij+zu7iVNFdO4H/YxBrnlntdP2z0oo//8
C47cfZBEQgvDk5qzZ94rFzek3xO2bOx8IrMQESG3m7sxtsNcxt+ePjo34HWZVOvOJ9ugzhCwlFKm
rsW3D/npvSSn7APMkS1kfi2kJsOM+X6krOjyL4brwaBL6ipmT6Fe5H+3LHE52znTatr8SQ/g8ffO
oOAvNd973E+EB41oNCECZ8uz6rdraNg07pFdQdtO6ybNeWRisT0tWEzyqTKF62I2P1HOWLktMH+7
DP3/esuFDTmExEAkk2YahxHFlA8SCotBABF9ctarti1ptMN8ScQFog7vSN1XvBHhnvZZK2gvOfpm
XRbj6R7hQGeE8+Re0Z3atDt6OuMxwMqL1MHHYNdpw9npwezG1bXOMsr/0FrMKeDTuCS/fvto0H9E
dYRnGokYoWgQhTpNJnisejf01UZza9W7FLJb+MOK75G3TkVT8JUgWfByKWI3yk75y5awQh9XlUAP
0UN4a5JdZ9CIRwWPdyQfIYMIAnbiOEokkEJcq2YDS0KYxRV4WmoFxlWVWAidiOUU4stLsrRD4W1A
Lem8u5WrvAR8ralN4SQZAnvUQh/pmkSycOwbBt2tgU6z6emhqunuvEMQL9gPmGzkL1HhnkVMaaJD
qI2n3oDcLyKV1I+VWJj6LCj4q1vWMJPnsHqs6TdH+QRLAyaxV/A2Us9/To87NK+btQMdLD2wnV1i
zLafNR7jTJvNVAFkZmiX7WNV3DoaxZ1qlAtGfg3EQWZI+ivTXKFR/pyAQkQ99sFxzJU3HPXF/LDJ
Y2RRieXyoQc4tU9HYPmkrC6aDKfNdDSjfEJBD5EsKzZotGbAvdj0z4a82PtoJCA5zWLxq/agoHbg
YicwSYTZNGcAZrWg3zWrUE1RlOiezw8OpVBMS0XQtvbf+x7quOuLoMJORi7qL4kKIXeRDvst7t2N
5XRzm52SddF74H6HIkiDM4KtqZp1yuGkY7hN1v9aW/ZTD8FV2UHZE8NnJWen8q+7rv23ICoGXAwh
Fnow4b3cD2o40RlK531JQ2OIIIkgQEWZBHt8tx7RUSWmir2FRUBPIlQWZSCiK/2CE4W60AfQ6xV3
4OzzSLAOoF73HsAzdFss5hCWelP/RD52SluHiQphhL3K/H3rTh6WvNCvcPKSfExiFl4ZuCHjgMY/
oTTlGQxbxkcJxO9KBPKY0POX3jecR969DOejx6BQ3YXOBFjiH44MhdRj2afmDfTgTJpJgMN+dpjz
t4ZJlo07ocCx8VsaF8jgflCiPjo5w1ADD+60vM6TD8YR4IYXx/OiE16/ylDFwVK7Fl93YISpVpAp
q2gnTZ/kV/WomBfVR01OyMw+iu2ZhG3DMjB/IxqW/l1lvZpffJW23CzgfArC2y9pb1UUk+VvUUmJ
AlPs1jBGMtrOugnzTtMdTSKvUpB169ASQPFa0YQnZVoUgZcABKGJJf2kUGlGnDPNE1PakXsolrjC
kKnnnl1F45+qZf97woDSkRACmg7UhYb09xfB8lkgh+xYYsnAKy8x2TSt89pNIZ2p10KAaoFKi/6Q
FCnQ2lyfpF7x3cDskAQXdXLlvXxYqEaPXayQ5NpaK9D6GdJE9o5sL/4pjnwk9dNa+OaoSaZ0yUux
85JT7GLu/Q5KpH8IwshK2QRCu0tQFvIXvxxlqJGG60ZDnG2MMlxD5hlfFnyNOIn9L6o2/Zb7IsW3
0TqheFbpX5fhH2uqwXCmLBU4sAFaIzLeIEx1NvhziV/2ESOmKKvzR436POTaTFe4GvlaI2CgKe1o
yRnwNQ9m+3pNJzTUHrP6veZ3IV/rdAEQU/zo6B/7aDbOJYKwltB9TFcn8Le412jKHcCwLqtUwbgX
8F9Oag7vLTIota/S6bIKzShq/SHFASnxf/s53zpSjzZaWb2r1MCObf9x1SldrRIYZPT0+4AIwwg0
vFGsSO43HIG8ZWDunNaOF/e1le3thrgLdpMACD6DVmNQIQpuuwPV7LJC46zV6AZEmzjpQrCY7Sve
E9+lPGYvwucZA/lciXFV2qUZMUAbJEuzfkj9V+Q4UfM341TEZm06Glyod5Jwokf3IbfU0POu5uc6
VzvBreJiD4ZYxANpqwUiz46Fis2U0mq5ANFmLhqbCG/BCeNFIJZJegdLYCVN3ptKlNTxAR6nn1GI
OvqAmHmsvbWjIFGRJX+1kDl3tk1tBjnQtC/2c6/ImCvFy53/Eb/lbkSHRiC6O0OjhQWVeS5+vgYx
x0Jrsp4hZq06pa9g1DKLdhMOjcdcQczJZK5VG6hAZyJzLrt1xUKDQQECxiFFR/2golMWtX8pvcuN
brkUNsSbIr8BvdAeYWaaX7qHbmBj1H+JkogmZUo7XFv3TSKaO2FnAHQ5dgMyfWhV5JGPw2Dn9jNo
PKLxKLjg99GNc+r/eWR64LplFewVxkwoICHMZhzwlH+NGkpMwfJ3Z92BwXFSqmMSNSeaJUfN8paj
O/NXouplfGy5Mj1bipxw7rYEydVDumnCQT9+U4ZGirkSQT20Uu6fsXR7VdfOqPPp9NFvmonD/cJR
GJS2SvrUPKSIhEKix6tDn/+mrlRqTc4PBiuuwVwAeQFGOhCFxLJ4FdbVDnxXsbjbsyLZ6OokUrIl
9k+p/DxTa6PpnaEFzaOwcVpi86yx+c42mwOTSJR1FXuDqbULFwmVJuTwBARmmmkZhuzymPSA7ZnV
skIc3zSbsEYAuejXgdpHIZUUU3pcEMrpwHUcbGuNvHNXfM68ee0rQgWqrAMeTibj7m/xKWN+SkZ0
Mg3diRU0AOUwVO5f0/60AiuNshxC1R5NFoA5cKKqXm5n66Uu071ysZ2jOx7jJS9QdhbxdqN/7DiZ
B151emk5Kg7+CE0J2Lk9LDcRLNiBNGeoEQ4N5Yyg4y3bxBWGdKtfkOljDpm5VdPkbMYt3babdXaD
t9jnW6gRL3BqK39LSk7i0AeMt866MPicPw5xoz97mHwRkDNdO4k1FeGY18ahN9psr7ufFZev8j1h
HdRRaxcAoqdObGSj0SY0jnf8JCndosb1+DLbb5Mk/EQLcpt8IOKjzYI7bcdAeIHG0l/hZaZtFxLS
bKj6pbgWgfIuxsvfdlOGJrrb0kLghhjWYYmFMhl/+poM1Jj0l/GfM5mTlIG15scikK0KygARv+PT
n/1CPagu8CZSBdCQ+idj1ONOgteYABl/Y9YZ4UFUd8Yktq7RPWrIlTb1eVXmHiuvk8LnDcp4COdZ
wiLknjaX/ZPLNfl9Phcr0YUwcMf0Czs+2GKU2f7EJSs75+6atJ6QqHdMbtIH3q2mkrsncWO2Bxx4
KtX+pLVpqZ0q6UTAJmvjf7OrCn04WlKtjgAuU//Fzvyd8gKDpIoFUpAYt/d7MMsSPsXI+Xjc9+Vj
hv20wCxvj6+HvuzjpyIoB1Ql4FImhFvbNCTcWg5/ihxmBqPzUuhOV5QPvPezrSUgD2bTzhrGy/ih
GRq990kdWlOG8FuvXe7xPr4L0cCmKfGVcyHzW2BLuAl4p6vwFbfy1cakOnTg4G3qGwmXr+SjRSut
WZLUcoJiw3Y6c6/433F2/Yd/HSSX3kLuHHj16H/aZ64reF7Gzw2FRW2YCkgyfH4OnGAMpjdufjcj
cMxDcpBX8D+2Dn7TzCetnvdST8mLjrf0+VBja3PyP3sVGEmeqYkfqbEcqjnDgs8BWtWEFWy9dyls
AePnSs3y/lD1f5mx5RtwrL7VorYwYgoxvknB1GiScsQlCzmkEwlBptEReHPvrPgrnHyGMTMW/aCw
ghbuQ8rRvopGwzu1OoG8fouVYQCi8+QdJwt8cDjH5Tg4qtW8hn4Mgbu69uQAmjNYlquDpE7/um0+
XUuS6Lfzj+ilX2acOYS0UYYwuQCYrOE2OekHgx7awXswJaGrYt8zwHtJIFiLDIVzOEbbI5LmIAY+
iJYQpeRq9eZN6+tITT4QfDhXtIMpFXU5A5ss3y/FWAkcZFKAw1rK91yoq8DQJqYZwPk3kpC+rwTF
SNU5j1qpKNaF1bGE6Ds/m2jUaNTXwAEoxRKjZVRN18XNI9SghYc1rauBKPQzkSvNvaTdpFsW0bzb
wwRfqB7pg5qFVz7t/RAZCM+O0/0cJvOhrOxQZ8sZ+PI7QWTpiXYl1CR3wBOrWUaH0DzOGBhBxwsf
WLNoyKL4mU19M26FB7ZugXVMVlvL4QycGYk3M6S7ZsFogqupxnn5tnX65nLoSK7pCaEGHPh8n2MM
LmeaxcW577CEVeBxVJ0eDTYEAnLHEtRwDaF187SbUK+h4dtGNDAElJVmcZ2MmHSVOP7AmUI91SKc
wtH/HMIli68QGPjBOy5oQEXjUWrhTb6rTlJXcvVXcoeCZGXmizMkpBvfJ70k7vNhC3/fIxsHA2WL
A636yKF7/0UVsvOI2fZE9zz1+cP52GL0HmaZgU1Wbb3HrG+5CCh9/GMmC8aQQqmhkycdt10MEU1H
Nft9VGaSsDL2WAW/g78shYpAOoM/uewVNV23rXZbwIizIFKYdsZCk5OTNo3yyvgYzme8X61W6l65
E9ZEzk67rydTbIVKosXNjyBr/ERtmlJ+oZgy6JTgBBGdYV5DMghbnb5Oe0EAJqLqj8YZ58Hp4oGo
Uo7AAW3jcS2tVS0MOKXJi8kjV2eIjptRuqnXuxNKn0CvXV23k0cTtWcUUpmqxF6hzLY+kyvBx/5r
PETN73NomBsg45pBd/j3K0OCdRKK9GV2ykXP9iLgjSHFL+Lp5RW2+kPvxCjOZrO1szOXsXvCgHbb
1VJutX7/FD+dlcczx53eR4WJfTi8X1iVpCIo3iVx6lnubFY0uUDAOWWE6b8cmY+5Q9HW26jOSxR2
s3ItCStVT3sYDpx0dPjseg5uQy7EuiBeuoOteHiDo9pXLhyyI3dCBZVhimVXJlKYY3XdFhSzpl8B
Xo6U3NvBaS6sm5iOwDys2PhnsTr/HlCFtKfFZ6qeG3rUwhpsHvgav3VaYsh88JqX472GHrIDRIpd
X1XaNUArpmluVQa7lXuQQHkUrwyhaD28rUGgF5n73NSuxZi3nkDF/97j9vIVOquQLh/1o0pvoNNk
/ClbgEwP28mvcPoJI+N/lWvdqyUO7IxVfoWlNaV3QiTrPP96cmYWregnR8NvOhQatCQvVfeXhO7z
kCyqauSNAUlVeH82A5tcYIAcPa5yG7fpVTIUNSVceJO/9PlnBBcBCyUOynWbvZvwSCLN4sehEdUH
1aLh6GQHhbBQLuruBc8K2Y4+hcrEmeKkr4hQG3Njfn1zsJUNK/+KiX6rTgfr0eaiPluW/VXGD28m
mQ7I0g2qUP5tUstjxhunslNZFq2CLuu/8sXSxoaZoqWJoHOITJrXu2iJaw6H3MMxE/9Q01bFKAfK
2sxCiO3Rqo49rH+nTUrh1h++pi6/Ie0GBUad6HXgG5JxWoyaPLIHujTvlEmEvSgLzZUx6X0Pu9nM
pevc1gq1TvMEDuanY+mwNBpLEjczpdzQuKyvWtRo457XSKUwOR+Nrs0PPwflh/I2A10yIqJTgzJj
VTCNOUFxx/x0QqNDtzUwZ8MiYYJAnFbVzn/aMi/nlnm3fQZPN0n238rUoC7WBVOJW9us4M4+b/3t
MwFpmIqbyKyYXsMn8L8Hgj0ucdugOwSzHcczdmgr2YyrzqZ73dya84AClKDtV+nXkHJYwwUBtSCl
f55Uf02x/RHt5ZMwYcYaV4NnVslQAv1cxxhFH6yVPPSgWMoytywc9+SxkYW1A4DLYrmdET+1I+vh
BTG/xiYhVelsbEMG9JQ+ZyBU3sCIibdwB+eobKXSuwTa1h8/ogzHIeZvCVr2ixjXcV9aPCHc7+If
Xzg8LHxXpwfaEQ/OSHjVnRnGON/tbW4AcyKLm1nZEt5h3rC/Ai17bN/zH7OMONL1QZzcLMSJv9zq
nloSVcIIXtjIt38lZgeFK9Ya9to8M+G8K7FusWoPx/Ie6avs5Bdyw0ytcXpajq5jYuMnXUDF1aG4
boyD6uvZS1Zu9xhLemhfpHReFO5C5ZGcjdx+CznJPPzZ9+ixuVOM0c7K1Es37E91TUIMWPRvZZAf
Y5EqdnsRya5tLkRuShbt+tYqxk//roedWubAYhMd+i67uA9B/Gf+lVB0kuhVUcIyfhzgpep6cLKi
rG4icyMeMqmN5aq589jLLDc2mGBzNXK1oPKAPxzKqkRVjAwM8yc6u7+BRafXVJLZ46vs/8M87vJY
6YjBvjZHh9I5zdbtK0AjEQiUn28ViD3a8Ey0xP3FLJ8Bb7Lth4cYmoXTBXvvEGIW+t7SU1caTUZ3
wj9iaUqvlmpIur04i8He6MQNALGlkFVJofZbhxFnYSb3j+Z6Lyz4bLsoqYKhk6ad7IMd9LxU3qtp
jmEre2fO7Zd62NSoMpJiKf35QnaPKdPP+XwF5Z8REchfYAxoysgRzRmmexDqECwAm7ISQVEDJsJL
cs2pKLX9HfKavrbEkYXPk3Tjlipf6HxHy8YpTpPeOvhygnr2nrEumkC915aPBypMs/s5Bv1K0GaX
n5IbtKmMMmIYcxFwzgVMNsBCV1YKhjToKlGtzGLc77HcBdQbmJyEu5O82QOyfL26dMH475Cv+aSe
T74rMxFR24BLn15/jeyuoBBRnf6bOEnWW5VOFvTGn9s+QXEFusTS5HviSS/QR3CXNRtBxvVWb+1a
xn36CguASXMWg73+/Us2Fpfp28YpP9X4oqjs5zK+BwbrjBxlgD5bf5lvvn7HuDRP7PtJYYHtak7y
sfvYwY+Lzg7umTVgK/4/CK3LX0xEIvUQLqEwb6IWW9cOo0+fkpy5R/jR6W8ktF5l6BjpzwzC+yhl
OIZkoQTWS87/MKU5w2E5kTYJdSbylW4+91lrMuNtPvPjnWK67WmrbwvdjrPUdznin6hIK5ewQUGy
nj5wt7b21TuGQFQdoMWw3LySeeSCFbQFy/x6WzDuw0BJKAfAAH4AkuIo6ViXhnSGeDspCYdhwRPf
JbqGpwWP43ve+F412dsFk8ELendRnowyI5VRQcBAuolH2k/Uz34CgEWvQO2CQotToT0XYOQ0fIif
yN9UcUc9B+Bli2m6CFaKwG7Q6h2T4NHs64RUMxCY3t9v2+pXamNDSlQxG0E+0ndlRVl/UY/a7LQj
n4jh1bqUbdM94jV58PVprZuBl1pdEFp5Zyb5US4Y/LdiUVQMDNdIJievrJcIB9+Bj+EJMd6Bi4BQ
UuOdofvw2rkQKNtplNL64GXqzvgbg8TLQ0vCXl/ut/Dw+ZetJtyBp6lraKtjb9lG+sHS1u0oAUK3
gnJENyhVTB0IpNbhuvNJdzFXIio/j5qBVSf2SyKODM9m8emW4uMEaUnePuoT2mUPQtSLgH2/v524
08fnWIkEoBMogTB1FibtB1Ym3vVEv9u0jDBDEjSqeZFXM58rtG0AOg2et/XDrpsFEXBR+kaQ4ZT8
bjQoaVogmQFc66nOoaualz4Y/5KtNAW2JUPB1s6gAEWcZB8XkENgZDNs5UX3kXejZcd/8R+Qa5AT
09SJo88OfUI6FT51m+XEiTE+UFTVbymupUf82AgkoR0IX/uPciJ2PNmAjno9HrAXjlEgPTUHnj3P
LwfCzvtJ61qBER329BAJ6QDZ3ONgQDPP1EScYwgIc1pB0xIo+KWoUTNLYoYvGm8bu7wD07rFjfhd
O1bdLgdYiJSSUZPXRU7+LYf3JOt+6j13O0G1LVJA+GlWM686hHhpKGgt7CF/vJpiHvPY8pKjks55
OqsWu3MDFLlHZYyyDCgz+7DgpHmS7I9eXmP11bZZMg0o0hsLZnLgj7aeeln2vJySFEZHPGYEEvSJ
+10DbagFhtveMVGLb1IT5Q8kwAzRqk1kBTFHCnsrCVW50pTaqrzKCWajUQFXneIyR3v3JjErn0oZ
HtiFE6hL3scW2qNqfS+aTrtysdlyFmtqyd80rf7AXbFv4C0Ml98bwZWWU0EXDBT69U0QlIr86+d4
DkwAp1HAK2mD57yIUUandjcYO/gaKsot2JE5OZhCmZNG7pkz+uu/HlO1V6uUfUWx39KBZT0MWaA0
Qxmt+3I9TFM2U5xMR5qg2ZTwIlyUz+pbovsNXdwYU3KXywL4dKYcDIsHIVYtN6OnZdvn9QI1iIFy
CgOBwqcp4hRRvHYwJxyXZk4YTiJ/7cTQF0mpx0Q5er6kVHib897Pzw72XS69mHaVidPJMyIebFy+
mKccX77IP9YM/miHdP3tMZisAO9U1ulMHQaXGOJmmsRseMWONEOS6/o9dxMXj2+VRl7x75kZu7Pa
5/vtvVtfseCr3T1UQmuTWNY7YmNd1CauXPQVCKuCnI5Z9y6ITDXqHb+Mi1vOAJxMILgu/Ow3bTe1
FgfKKOqqLf8b+Zcxr8bVFe9JDRevOBJ8Z2sSXb0ADYF6zomgNZRVedNRFdsx2pY3GeV1TKPzrYc/
tpKpgBkx89611/yb1V0U5UReXEldyixBBfr40THxEgkAAT/cBgCnYoBEhfl/BT/vBndbUm33YmHx
bKlGlvI339dv52hw9uZhFVQtQZ3UadGKb8YddGFqzSOpDY7yc/oJuZB6qYQKK63U3Oaz+zj/Pd9a
/tFqTlDTHTQnZk4+L+smlqqk7JOV0b64iqKsXv5ve/JoudpTFUsqmD5aciQi+s1j7NScsfNierCX
6HWgXgrMKcIji7jouqovUPVUCQfpvmyB3IFWM74/7mLuaqfCrVlyadiQuJt4jaQ16xL5qEpBPYry
foMsXgrNEDcTa7ITCHLGh3PUiG4ol9mGGUZB8L8dTTa2ttLpDeQLRTjdoheyT9lOflE4LqNZwH4t
uRTwV+iluArY3p5T3ho4SsM1DpFjZduetC7zY7pn7hOY/UnjwIB43mFgy6RPRU0+6ypw6w7P8oN5
Lou2WPJ+IFpwylph9rUtxKhddcLY9rgWUv7ptjvOM1Zi/FYXCP0+Uf+G9+SoP6Kv8hah/YTpCfwx
9UQH6qzJxxKsvLAxhyd/5HxYYoaj5VLyb3AXbbzfg/b3S399PJMWsJOMlsrcNxN7W1jdFxsN3lop
f7uywDwpKRSALsjybUvN+0fNRTxshW0eVe6XNIIPps/YR99qayp/v/DuZxnA1+ZyOzr7onUOmMSy
ggA/XQc0UXCPDjlXxt3a3p8sBlTwgHDnrJjZR9VPWvF4HKZqRQ6b9IDFOamp6WfAnk4/1fGTNitr
40Kx8TPfBWVqUlfVbDrf0jHaTBF0izZwnN0Jrs4bFPXPfP7X08ev4ArAkJDNamA4jCYXbKe2a9pD
9lGMiTeWsbAEy3D9QkGp/c7AV6DJsiAIj7s8dPH6qJ9aPCXChw+zXSi4/jiBKY8mzQa9FIgnENgA
FovkxYQQTKBgw7lMlhd5qwIjCOGCpZZeV4KezrJe2kk4CcuJACZHrbGVdji5fsQsiejE1dNFVYJV
wpcU2ASRz/pVByAJOAktBiOnTkBzCA3tloz6RsOZ0arrIgboVM8aDNjF3E5mefUZeKa+26VbAJkj
nYD9GyRbTN2O0aDHb9LTTjiNe8BFYxh+uP3ChDnEQNfRvJEc8pR9+y/g2c+AOFDH0XWH/T7++D/E
S2m161nKXoe11F591BL0WDWDXEbqqFPqgv2mGuUWAEzxa4P6i/POPlLflyZZraBdzRMr1e/B3bjU
E6Js24l/tyIEHg4GmO8qkrU8gXwtOuZdpLrc2kFwkTE5fSuQBykWezSQv1Dr0HqiBHFaWgOWSqN+
DwhQ3P47n1eKIfkXe85XS1nlT3b4cmHC2c4AO5Lhc/ojCgsanmN72XS9ZVi81k1M1XWs5qSfBsX2
wgssFGK3lSzMsugz5rzEQKHH4zFLfMd50H0dgcCiQUYaGXl5a0PAQ+3RY4mlolzE7rAFlozS5iUF
rjTQiwzgiQqVT0Tm3ivP+JSMLbqPLe8nyrAt/BPmjZxtx4CLbK58h9Fs1P4ZwBoVnkOTtmAxk7cK
LhSCbka41IMThE5/Fi06ufWJ1XWNl+YWZJp8pPxAI73E/+GWxhepmWJ+y9mQSkNFLb86dzqTA0q9
I+qDd8LCgSUq2JxEp3koq75ejpKCKO3BPgFX7p1Fl5fmilEE55Oxa2ZqsLuhEmZdch19Y3hQA6D3
I5y1TYb186Mz/izRDAC2s/L1oSvpG+aCikHyvO5UhvtW6ff9QPpuiZKx5Rzz6Nz8EaAyhQc7/a0w
M2jf8qZ7MTPYVJ50YacNIRSNB/+pL1WessDlJKayGY/xQrWYUI3QqkXYPloHK6lrfmplnuDR3BhQ
4KiusS2w+z/qlc9DftgrjSkHR8fwsBriFjZt519g0VI4qtUIWqVTwm0RvKGpaj8tt4WhkqCQjnkw
RhjMcrqoYNgVXeHc2J0fb4tWwytmzVAiYTIO0pDkzr6zAXkcE1GC+fDZ3ywmKd5FvLDdl1xDeiQB
L7f63MY58zWetWyWzguRg4+NP/LxBonpdqugRB4ywm4ZQtfvjc03a65HnGAJ6WEIF/bvQod0LzK9
dwD1ZevXGxqM8Oan4GLd6H7x/yP4trQwLzJSUbhjCvw6/ln8Ssm+WRzGB3O2kqf4y7y12Vn6FXtd
Na7575c5WRqDhvF657SuQHCqgdVj/2GnSPH3lQY+dEBidn9zJ59sUghUY+QJ0qw2immT3q0EjKZj
x1jBIMbVE6CbeeNH8Bu791n6UvuPrRpqQFwo5ymLPM7Mg2dt9Bg8CoTNDwnicB43SakL9g/sQyq1
spmv7J6aSd/E26tqVIADp9/AaLSCsAmqAmOKB+7tcKompWq6wndbmzY5iYXfbYXwmcwWHv6IakB9
pxqFjJirHgBgLR68DQjSuGTruYho5aMj/zRTklgEUscCOp++uAzN8OaaSIqOyvixexaPy1zmso6R
PT00DPKAHzMAh3v1+tr6QGCnl9WLhFtD6rml6w1MK8KZL1l0psryuXtssWjwNtbGwnAOxnXSPX/i
5TFbAADlgtEfn2kCh0LFfsgh48548Re3E2QoW2wpStc2UBh2M+v9i2v0/DuRl2vY390nhqQOkh+j
dMFUjc+Yw/Z9sW84Xs/Rn5z660TWbRoMVc8ny3uu3z384LGnbCmL4+NtslHu2LNZfLgUjX2wI/lq
+wRajnKzI2lDCa67TmlUii3z9bwkdJjtedJphOm2MouXayIsYS1gBXesNSfQCN10zYDl97QsO/K6
lFiOpI7S5y9RSl2P0zLbfECyx1xOZBQHDUuYBAd+spetz7kbFX1PeuTggJRa/UYeq2I+ab0e5ihT
swQQ7Y+BZod075dWA04JVgoCs4MmhP1qs5HeOEs5izpjiKGgESux/sn9LJjRMcIVZ3lyNquUHNPQ
e8bp8zYQKBflerM4oFs/i2wobF+OrdJoio6fRcA+JrvL5h+ymM79zgAmLcT60peuaeRgd7dSvfJQ
ZN9mMUEV8PHmof9j5cctTTgmvVVDQtBrKIoz3f/qnWtBVK3jQEQQ3ok2WxKZoa+ztRsMJ59RgO5o
hraKiHKgFuyG8fKsRkpIB7GadVZFdZ6zoVYwF5Am/j9TbJv7XA7D+diwHj+dhJMELO0PhnN8EKPa
OLIGShYVQbtqDR7irWk4OnB1ZpHmf1iDqtwS9faTgRKnugKFSA3HQGYpog6c1mX0M4jS/RJ+Vk2v
oboknDrxNGVpZgiUJibJSarjGKmO4HsV8SERJBj2wkK7EeRYe4WyzgcvJxPlY1yzNJgsV3E8j6mO
K2ygi1/4hwG7MmzgIgBf76vnmNOnDk9/tM+aEYCLR+aVLjQUBgk/5fssNdmAluZ6QTbh3IxzJmf/
AD8ougmH/wEB02pBYr5VYmvHetDACMMFzv1T6QC+NAYA+3AKejKFqHpg8dr85MErnKG7leT7UzuV
pMDBPrQ0fB8hvfqBEmcZcG4Q0eemXDyqQKAt0jOSX/CbH+hcrnxVRd2DdGkrU1R03HLmDn/fqACo
R1cVkCxeu9xwGAy5AVFGguPJ6fTpsyyXhAvF7srdErYjt8lpENZ4seQsI3pBPhiXWKyo/6IKicwU
SyI5pnqnXkuyhremBGUIGa4Ft/J01upQYrWfcyN1NnXIGA01aWZmD+52LB0rLfyqZcRT222FHUJu
NBcRLfEY0MfpyGyx+S60+si//o75MuAxvfG0Tes4EckWjJFq4GELgST7VW82s/Tvh96/TRDw5Thv
TM+y9Rd7Kw/lvr2kyN7JN3E0EkdvVtunZo9V7n7UkmXibjgRxhwwtlCi8SFarsUYSK/TO+FCrxl0
3K/0ZEmE1+WKKifpUeFNu4I298ocyQbXEVug1/AgUDe62TujGKeLrnpbb86+/a6NaZeRweq14QKE
DqrsqE4nI3XjhDF0v03TuS4SQBLWr+yrjYwUkf/jxBmf8sHThiB+nVSQSbbsZegRHaNZgGiHByR4
o+59ONn1NQFNZrqvBvBzE6h5PTpBe3rsbGnW2ZLQxJtcQJstnm6gjvZ3KP7b1gL2GZpLTTosMTPb
N8WWU9lPOEtSPKdG5aUjmgBFoA/X7dOf6VMenkePzcwCVpCfrbRgPqSY1iNpK/OVcpI7JA2opE4N
SEMjo644qZgMhI9KxVPQeZscg8arGXdcmaxyuOyCeXZfwjYak7hZFVK7s/h4Elx4rnO24tmcPwy8
ceZl6x5PT/ADKzZQ08xOWluXj9dBU2uyyN7VQ8uKVUPRl5Do6S9PtYDNfjiSjCNF9avZCKspNeAY
wsvtXg9esYoth0fJtJQSzUyWh7da/wIXz9YZtNrUP0g2yEQOhzGG8Cf2GkOb0jb2apyY/1VNRxD8
L2Z0nxOY+MilegwRn+DbJV3Z5bp6Yg3hsmKFVIurMRDLNcwfTgjqK2uKxK6rkXX6aCW/0xELNQwf
ytTU/rA5SejhGyzEFz8IY3Z6kDrjynT6Yy0NqOPuaxQIYJ4On0PBw4qiprptVucmSScL13Q2yl8z
E1rKC0wKm65/AJKs07zwBunxl/hT4SAiOYpNKEvsePDoS8PyYAdy4FUGz9vykAF1ceYpdMZdtiNe
IDGhyStGdXGNy1hLnAn5j+fM0hAryToijb/lfPvdmorIcF/908JT4tQkL6+w/jGpu10glUSmn12J
3SPuin8B5lEZ6C38YpW4r+IqUUZ1biNNzjlgsHzP9clzwjbnlr9t5XATB5VJQDwUqjBvDudqzws6
wMi8zL1LGgMP9me/s9a1RVYARAvSPwxT1yRkJAOawzQi+8Fo0Fe/KECThXdvFj4IIHN6mM1tLMgs
/UeIe7AIHI0DTuOeoK85gYRpw0WZV9GGbusQbcd5kIQvby7k8Vc33xbX1nYTRsVbckgNPyf8XJ2r
JgXMDOKNhTA5SCJLi1zf7z7i8lSjI3nDN+5g7KF0jx3e5z1US0KK3RCbHhs6ppHN3nj6bXfocPXs
joH+TWWwN94sR6hH6NRFJwCjoEIkHdha+xIZzZxXGzl0PoHYWEpk+rQ0JBe6Hjbo+ga1FjFvqy0D
6n4HqalzqXkB/QikQS7Qcj7xa9OmcClKu6RvEiwGqxgfLQFxfOgKOLqGIet6WFOYWHeK+6Nxvi+X
nP9Pa4GsX2H1RmddNfS/uF9YiLp8OmYzQgCLUW6lW0vLLzc2HymvX0qQ8fJJk6u5mQf4kJl7+Mib
8cqffEUWb74yBDwOk0HvDiojZQJ0MlLvfNEs1KT7t40QuKEWAxMrcBPuFiE5Ue8O8rOvW0/6lPbW
wjwoikgYMQXMB75TsObrXIrEdWDbRkrIuEhAVEB4C/grKHm6TlzHb5v6mdALsH4JZ06fZMZpUmI5
+fiGgcdwCWzgqbU5ZjFWrOe/3IaMOznh5nNLYHQ9qlh4x73y0V+PEUliPgGqsSyNE1rCXgEQ4AEv
boIdqzNzf2RSrgXMMnoRBXjlXHSrKPa/OHuyN5T4J9BWbeb45DFjTs40bw1a2yRc0cctZpbZKBu1
gDHG5+wh9rC9GAZrru862LI0HnDASQvLJcyO9v5Ne1dP7u6tyJX460MaFf68FsszIONYe7LwcWVj
lFYQ8yQbGlzJWMUepRbNdY4hnRyIkAs0RfivkxwY2zI3s4WisHHdcWRQBfRCLXmdIgeYQ62iOA1N
4UXa2x7G481qClHqLk4rE4Ix2V347ZJ8FGt0RJ9cVTr0F2Mck8pWxDICkbW8Hxo32pXSKMZWfsFL
RhnSP0ufC3wHJVpq591PpJPxG+Z1ONw56yEYRIHGaw0dlvHIW19Yg/pk/trzmwr9jhGiuVTcZi8z
jFYfRm01Iu8IgGNsH4air7TWEaNcoKYwQl/ykGdaP24T7dhfzyqIisuozclinP+os/gguztasA3E
aNhWsjk8T7NPceys+818OxE1bArF3NjFQVK/UqMlPppH2nucOuqoAQ5+6Z3SK4WeLurqmFp/2+t9
AbzJBXZ1yKj+dlJsiUOeVG8G+RPn9BIhqDsD84IOp5/153kk8Rysd1ZdnQljmr1in9RYMGvFzfi/
G9urW/CYiQo8t6TERvSzgrmGlGY0prFBwNJr6uvTL41Y5dgEezQH/rYBUkJWvYsdok6/onZqEmYf
9ElJHAjmSRvQa0UU6BIAgj66CNXj7hXgn7hZ2Kgow+/Y/T8itvqdPd90/1pJizi/ZGvEotB9PZm4
lhvyRmxmRUcyTzw37ybAs3pzIZgfIl9ECaPrHHJ+SXFbUJT8Z2g2iiwV+i+VtBMfqEs5CHXLDzRM
rrHLMZGvW8rk8iXJ65jZHJfBckmc1dvNNRG+8xDJI2vUG3mya0jbUngKPKEzc6WR4cCjvXfiw3mg
rw/P0ugJvZgVCkziXQpV50wOPt89TUwaZs6q/6Qxd0FZH7iNQSaa+IrsKK0RNv35QYk3ZgnC/MNE
VRA/2wRnreSoQ/IYTeT1IfteZ4ROP1MNA+jUXth4oEFvPyf4FXPFJUm4bmfLQiGvUI76NSsWeiZt
cAKOr7wE4AJIp4yXkved37F5hA02OKWPQU4h93o/lHXTelqqFXGiaZITPyvdQHdERUQfK+4Bhmsp
xPrXhmbpo3bpX1V2+454IwEJnIF8Y4y45O14srXi2yV5ZOsShzhgTlLIDDgud6904OGMhshe9VHR
CVoXt5xGMJTR6Wt865aWvsnVSDSoRTMiaJu4CJwiHhK31XIjsVvBCnPHVPigsXthUVjG956Hoa5o
Jk8Y/8QWKihr2J0WSvPLTfPBp8mJXfd7FDUn73OcPwVPqAcwkw94x2fw+/LQzYxTIU460wN3Lm72
q4PO3axB6LEoUDZ6N7OPjEfmGho/SXTTgFG9a1WSwhuPjVdZyRZJQvhsIw1elHAlhFqciT/aEzde
KkKrbqQ9//oaBsHBFcuqXyjo8eiFiDVrfco37ibS4Xn0tVUWRmd56psYhqrmEAr1urmkc3OXx1sG
DAeTPGLuHGcklY8U/h+GG7QYARjqG2EjYLdcDLU/BxE8Yaakkk6fTQ/oP8anRJZ5xDJx3AtYJshm
QxeuLSSucPNjdoqUMznXP/CcGAx1Ie3Flnx1Nn7GPRLdDSHbWS3e7yPFXuGNNMbO4CaffpJp3ZYe
mTGU69RQzy3PvF3FRNupC0KsvExM+BpCL4t0Z5IqWBPOCyrPDYM6iBK9QKiokYpBMFX7RiW1C9ok
+QmDGEvy+NGpc3h8TPt5kVXT4myyANW2Ta6rGpJ9HJ1sdLiERNaD0DR1KiPZvmHa/mg5LcRydsY0
70d52xpeD1B+AfofhYplzKZfMRXtwI6MJl+kn4rKTKhN0HsDNoer+hGCf/ZWEfBQyCyltEMVAbHQ
bmH+mMMXHCI9e/KSoT7huwLlFI3rQKf7Up/f/wtm6dIcL2ELjeaR2PO+BqZ0nEIsLv7b5RlntoLY
8miOgWWe0nF77yhhwqcS41sSBQW/zk7/+M+1vsA60iBKgNKUtc/bVJkdvxi3+m6TmY1v/nmBF0h+
D3cFp+zbPXMF+Wr4WBjReICKW9LIcLjLk4cGl2AmmdpeNZ1U+uTHWNggM5CmyAbrM+0jz9D51K34
8ye7W08rfEs/s3hXaqbQkAuMzQhQMg9qGZgkPIyXz4J+ZWbrq0LV5opeMCXNXVN46LevjOdi277y
TWq8I9nCcBKkf2rbcVu8vGEPJ2LzQfrOsCxVrwXaccDxA/O41GQ9hT0cJ+MpjjdbJ/nojPZWFpg/
L/M1lZAOExbJe6+bRZs8BD7yLol9RaUqig3c3rfiVkPs/DmnvawxrbKpLnsbr7BldWYuMnKPmShd
FicKxbY6jpGh6SJikvWsyidTID9JHZC3Cg2C0qKL9aJxxu59nY4h+q0rAGteqLqoMjkWluL+rGva
dPl/YfE71dg+tpNECVGUa4SjX2qnRlkJ2n08SvdV1O9SnQwucIWGls30hP/mSYoNifn3zowOleUK
PlVU9p08McqviFBYSEagnPIZ0gum6cYCNRhOOBzOHkreLvTrzamxfR82eMglz52/UwnwlV90ZZ7X
uw19OaZtAVKEJE7Tp43c6F0ywcT/rGN64MbJkY7QCKnz9tduZZaJ82bqWU40zDpDeXysJj5DaUN3
JuUpcoU8tDaeNEL5KLuh0iGKhYLU7alAI0de+MVp3nDsXPDz7/S5FyXwIPCD8DylXrDrfBaFDdq3
FkF2iGWXwt/+wr4Tq7mgt9poizGKZyBvwKYZK4w9arJ9Dpl7v/NHC/eR/zEu7PRjGEsnlXSYT/8F
6byMDZEODaSIByHyD9O83FPcv3gwgWK+ss7/p4c+POju1cSokdKUWuxK0Ok0dZGHBR2YXYnRr5EP
MbGwM9qL3kOSDKlUX05wNtHYzzH6ctKIA8o6WyiM17sj0RShv5CmdF2d9/Fjok5t2HOGGF7w6BFm
ZyyvKCWgPBhImC5jdGw+L1cQy/Vfagjcv8Rp/RfjrowvumdP+tzHNbnAd9CK+Y6d/qDIco9p9P0z
4n7JLy7ThGn9fOOi/55UWhlK3Qehqr8JpgxKbO470iAijx9AvRnCUKF3tB7tQ1AGz1oMIlcSSgyt
GfVFJiYIWTy0IkblNIM17B2SSywIAHRT1DiT6TsJsWFM2uQqcVG0ByIHaJox2rFpFayTTH2dCQ59
Txg5ogffm1RuWBefZqPnfTFX+LkFUwrxUJDJ/0I0UrF71cmGvUe5Qeckwp8wwAdWffDMT/TMp04i
11haO2T7qUksiS0jkOAkwk2GIISdBgGfTzyR5TiRrwVOPP6hZ7CXI8G5Rb7O2X+mj10eFNQQ5Grd
9P53frGKmRnWqJ1Pwv4qJoAvvRgCJoK3nIwKyuweDSOhiBXv97QDuimk9L4St+1nnvjfqs6kzK2r
iRpsFpoTNI4gEuVIRpe/MfHikaeEgaRFiW950mhhDjKlZaB0SFa7IU+RyRF92QyY2HP+n1AvCC/q
HKzg1CL11Dt/ZI6PQIPrLHV51bcg3Yx4RoNFlLg7N04+7sSDGOH5H36YXzwIAtsIPiqeTOLcNpVy
xU6PCltaliupdfYhGVCZp9oiwPynAJ0NTrGxa3PTbQKgTju5VGUufaWAcXzRco7dEh4ZPlGj+2Mx
eiVg3YGIwFPnr5rVjYP/1mLAXIL2Xc2uNN3CRJuMcYejn+efL08Sfb7WeiI0x87eB49furZdLQAx
uDa+qOyQMFaqzd+4Mej2ylIr7eRslmA+SDn8R32JDHVLLf2YQiEIwN5yBwLfiJUlQ/dcQvfuQ/o+
XYM3HktDcnTmPJP9DEs8p7uKTUMNLPMOwxEVr7A/J2jdvfq8A7fVin39AwUTxJVLq1l2/jC6DCK1
tsiXokuxdtriwWyg1w00P/6zO2J6LhST8xFv01CdjfqL9rAtbLjhlHrgzD4Q5aK4TABfpjzKv9n/
rop3eWGoSESfzAOZPLY59n7eVKALAMKmBE1IpYZpovgN2kh/tZGPOqe6KmWZ5TRAd61sWwSbLjRg
P9bP7r2aBItbHdrYgsndSw9jke5KhVN7J/rh81cgQ2MaSUCe6iuHoS57PTO4p9lvODghHeGXLs3N
lSHMXomrUEbJWnCXdJr+VRp/6PRTKg1EP+cxawJHcwpqlBTkn3ctZAP+NX6v8UtdlWBmkFf1DpFv
lJVs2m9eFt+2Rdo96DUM12VTlY4tUxbr1LVllNGsvVJi3nRkiyUhiwdaFSFOwo9og/7JVvFk85Wg
ATfIqw+8IYnLbSP8Zla3T+H+ByQTA8SGrL0urUqIWu/KHsLn1yG9Qezg0b36AHkOa5CRQSL+xkIW
3E3Ook1H2Ik2IsxMY5O2rXzYpOlD9/Q4NaG2h3zniDyV17EtuhD89p8gZeff6KXRJ8A2OnP0Z5ee
IiKodQHn9s7hzkWrRt0ZYY27vGiQPWIPxr8MWrQ9KPIbXvVARPr52U5/GZYrR/uUu4mWJBCGNAoq
7KxGjR4/cPh8ZmagU6AtrPco1Y7FbS8/0FlAgsKL/4hEdICxulDTTNe9feWSrCeWIGWjow1T/eYS
Orq7zqpA6v/mVM7Ah968mGXlusXejffbtI0++Q3opktx4TDK/q8wUpRNEIaNKwbjt1HAvAlTgPL9
OoQoNg5acQjjghGDwPbFi+Vxx1HXZAqCpNWADPFnPGTXC3SOPSlBHGdqEaPbEfpQ/kVcB8pOhndJ
1Cg8MBPFaw7fOS1nIOpfIzsFuvGGNmwGgmRbCegYHXM53Olk8xTPgd/SYFW/KiAKyfTGL7kII2tV
vceoWzvBc0SLPG2clB+R+ZeR+sxftmnDkwYEOG7VFGqIIFbdpp6kNOAVmFb3DhgenxDyJKc1k5X+
qFpf7Ss/JjGiU85zysVZJm6x1J0dOd2+kCKudHQ+/zjnsRryEl8bycwk01MhOe1Yo/Li7IQjCOrd
WR3kNRda/1QXAmMshhgYs3ADLak16tqu1wFrs8zcdeevkKS0yyKzGlXZPjVU1BApMb//vOpHXt5Q
76zNtemq7zaS795K9sOoMUZC57YPASQlcop0KCCwtrtx0iIK0peA4HmuIGzzqv+iwjVfKhviiRAI
w1CHCxGSl9M11vPiMN9h+VD0N1iFx4dKuEJC5CwZFU99Uq0GfhVvEWTfDomAIHbcRZk8XxP0upOV
l4Ci8J9wHl26EOc599u5c8ZPtpnJKeoWb9rI1LRkhYtfn0UypLp9PPFIbRn4AQdGE0oaR8ErLm5m
Hyxwqrj0LKXgFKN3xPR8cRaDEPRse62AlhMOPULGaDlV8D1neyDk4lOGPYj81ofOcpwo/ktgr9Gv
a3rnRjzI0RiLALXCzmh9lamPLZmaQg3zOqo4pJ1XdYOiBy+ik7AxgYmob5YTBdcKMHlEA6RqwVw8
l136SZSbrTJnSJDpt0Y3a3jSXTq1Jjqs7UxZ9pMSBOiCyJ+F4KLoTmDbFpbj8ruVrdFQgTvUgXb/
MXlZO2zykzMEqJE+2MR8q/dvopjIWYhfp/MHtw1nX8tbR1BL95+SrCBTnva6Hi9JiTeL89CI5441
Imq1cFEZB/4xgZH/QtLJSTctsaYvukSR5Qyap/EDmO4TPsViIwGzm9DwVr6e4Op4tNpry7YHjiHP
xTu3/DqTzTAj6iszQba/fFlLz09Oa6/7OqJ8dxdYwzhzH96EZE5PEQJL++UhAQKsfWINVcrf967P
cOrz4Pyg9tKQwdiAlKJWwdNUcwo3m9sj1yzrV9sOwy9TlsbwmWDhppFd07BXGJpddSDY2KZnc5B1
Ns8GsI7lAnOfyt7ako514kzNHR5XvxEgbcleWwYz34OPuUqXcQmwSw251Xb8/PkzO15BqdKXSlhE
KOx7ywJzXvODk5Rp3cXWe+PZVBSodE2aEXkq+bc9sfFxqAAhfqZDmbtOQvVK+t5HAan6Ewq4yheM
S+OOmR+uv6ObBJvTIc7u6lY/D6VrOYr8zabu2BkF1Vh/Yhz0Q6PC5aEaCux9J7q1BrXRySqpVXKf
YJmEatGhnI5pt+b1Mtssj+wL+smATsSOZ50UjJHPGFpP1MWmV38ItfFPLUyKar+dUQQg4rbRDMs6
BeXcz4E+zZyDXeXkl/Tf9bHPNSVTkW6fuQq2xzQbkJy46KDnj/rirRhrK6pH8TR38euHocZPTu7O
kpPJvNH7kkdD7gJjfV4cbAWXHIZDnEuiA+Ps5hM/ILwyELqapp3XCyPjiGbuBDhxZyqsnzgTgh0T
xeO5fV41Q+Z/t+SNkcZ7kX+yNjacfrE6d+ag87nSGbayuajSgqLq84ysbMNdUV23diontCT1Kzin
d25C3veThTQUjwXprbZu/ia/ZsAwZ8IchJGd54sACccxqyBeyECj1qJ6L9ovLYYm42sB5Oxta0RE
eiwD50qq15qKaqUDlrMChJUFlppAQ7YK4a978HiwOR8CF0NCsM8z1SbbVshF2uhy5CR93ibvUxwx
o7Kdie3ErZgX0f7NHYD7PHCmw/qnoboJt9cVjAlhRjDmRyFxYdKUpYm3JqM21m9cVU6bXmap+9QV
utdfE8vXnoktNyx1NmAg4g7CQq6bqGrw3CvvhrbZROr0DM0VNZ23aiyRwCxMq6Z9yY3bEqJLThye
YzUjlnKPWg/vyVgQqr13HpnKwB3avOpAnM8gCqi5Sk2IzGB9e4QQPsVxI+pphpVJZIh9OL8JoVnn
ujCOz20TqfdfvLlHy+E31roIMebxdm8JbsMC4t+VG5PTBoFyxONfGLJm6vllGepmlgLl0XvFK40B
l2CRT4VuUBaNjLXMm+tNmx7pBeRD/MV3P/yBxVc0wXVEBOF1bD9dLH+fSQsDuRc+8brXZtJIz5gg
EdTl/GF8NYxCVrBD84C1BhfjOMCa8fRoZCw+SwW7W3i84exT3fI/e06lo2REzSAeEVJ2035jqM3s
VlOxceno6V4olFAEpaZSzA0IubKstVHhoNUBgf3ebqYmXSIFW5vhJa47dihYnNCpWCQlrl6v/0YI
QRtMZlH5QdrV80Kp2rg35GKQiDPF13wcXq5Z7fXtl/d94bQj49vOF22/qGzSgeOpJcBZ0AsJGsNe
P7J5ioTMW7tKL9ds1YyKFSSFVMWQSMwnDNXc1KtdQ+T7m9lfaHEd11x9TwxE2XzhThQny9xjYJZO
zVtkILAWAUmNBNE+KFnqqnKO3ShUuSgvOgVnYwwMg97fcCpByiGWRG27Hq5tb3Sh2E2g8r8nfyto
g3wLeCnTWyElsxwlbMTBzaBeXtB1hKZufYzJoMYQur0BDLUB/zTFspOn2LLpYDFHJi8VbWh2fBV1
wuRXZcNoYQqM+n321dblOdzZpOU5++o9jLmaWmLJeMKmCFCw8+tJNW8NObqKeOKvyUiaddCXp0Ic
yCMMBfie+YJKya6kz01OF0gi1OE24BG5wHjzZfb6X4124Z4dOx0A+1Jm3E5/AHZ92bwFZj+FKCSB
Sx5ICBGQ7/9yRLFbQMt/PcrcrVdhXITULYerkCB0pa8XyEBk18aohlMlnpfiSZyF0omK9YpSVyTB
T/u+7J7iGxI5t6qNWHiQ5X5/Gp8jAUAikEjeSaXrb+WmiN2gP5hLTscA61QqjOExAIxU+XRYrJqa
pGepbl+D/9ZsBlE2vo8OM6wolHYkU+FmXCbBySl2zAomKOWm8KNM+TFqaX77kMIfiDgmi8BCCHQq
8CFOdXPioAA9iJKn5+UfzVDd8j4+sdd5lvaZj/hoCZz/HghFf4CrXM+9dJimRtc4ZGjwsDIaEqU0
5iiNWgf1ReTUYow3KDtUb6ORvXGoCHIxgY1zl0ZN9G39GXbzkv2EiyLknq7FrhO28ssU4Cj5+ZM5
aoKHffMsSUbZQ5ufcO9POFzNBfUMjvDW+OWPjXBZVU5zFuTQq0btqU1LL3Nn09n7uRH/fso9TKmK
FCnOCY4UjuiwTzncAwRvI+q8LIBspS9EudVmnE/dGKO2oLNklgtLx/DgopIKnY3wxaihrqEJljOH
uwIE7JdlakDA6/NtMN0QkEexdCmSkvz2ElotbKaNLHiwNozFheqFSCXJXquNmuLjGFOqyYjyJjDY
MoMHv4srsoHA0PHRJFqFiHW9xX4d3/XgLTVtQ8Ez5l0gN64fQNzdorbqpv1XYxccDIdY4hRx/jAU
2yZA1mQjibMk2RPiepcSkMu8ge7UWqlekycFBIzQXHR5aEBpgIFfQAxE1f/KKvzCM+Dn1F4cmGy3
KwYX7f6k7pD8JQ8BaPCh0N4R0ruiBlPrbtV9lKVBSbicEEY8gB0m22aWPj/LFHNwni8OVyMaWvhe
QL2WHy79REp7JO89ng0qm5/BivNPSdzqYCU9NIr5EdXcp51cqkeDNFPGDcWgSO8QijtGNCeEzaxu
CBu6m/tJOK+cgyKXAhiRMwIOOQ5tktioxriyP/UJNChOVLmLs1/08KdvQHNwNUqYdvd65w4IXefb
pqLYUl/9sH5sCOCvzJiRVbf2DflcauTiOY8KGh57tQD2Fhz6dwbHavoucUbZoVs32IeWE1hNN8hs
lmjzJLF4F44ko6CIE66RGgCHWzT8eE05bfP8vWlg7eucbM/r/8IcOUCm65LbbGTuciKJfanumZXO
+QmceEM2Tf/41EM2dC2FR+aham3Ck42EOtZkPdLUJsbs4MpJe4Km3y+RVAbFXIPr89JtnyzmSUvB
ib8hyimbFJhbCoElvZkKTLCSxd6e0C3ayOYbT15tBYhKrgSQTBugqc6ng1ye9cAKiV59NC5cUTt0
CgOrg+FJ93eZkmJwBlCfpz/clnj7d4hfAgvkVIWt2TPmgBFyibse6dbY84x6KiHIvfslOZsSBUa9
dqWFb37W8MiZdc6JgLYfv3kyvcPjlzxsnXsMnGfZ7cWqvJ6qyP2lAVmqAIneBhUCVjAXheIX+O7e
Neb28VzWYY15/hj+GkKP+sSmFaT1AFsfaVMNyQjzUG+SJFWUDrPOLo8bt6yvSJNCQ2sqI6HliWKZ
4rTKZ8Y0BgbcX0KEOHa/ZZa+VqazQ9Bz5wBCA9EFhHjhxBNBELxIMJY8hGt1anhcV7Ox46JkPULI
TvPFYPQ2haGycRzxRlvl2YGLBBSnTy8R+wkh0k04HNr9lQvDsYf7CEEQu/IAJHX7zUQy3GgAK1PR
WU/2ZvFBjq6NCuSPSu+4eTj4BL8Z/HqsbBmmlLgOUJ0LUkuliJ6UJxGIGAyNpp9RXRAGN7PeoO7Q
dJkv7KqIXegIwOdPTyeaODZuSGX0Qh41XWxOFGYLRuaaEzT1etAd1xRVj/k4vSeLmSDutNNLcy/r
NvTw1LkvfuLgMPWZom55+6vwzUDOTRr0PkpMCxxUjcnnBSk6Ln/D50Inee9YaPd7fV4QSX6uLSgw
GHuA6eWQJpPZniCH0o4PqPoX5Z/WN2kOwkL5uRnSxeAXIIbdrWyBYWRraMJNZUcVUfqb1W39kQ3r
F8IMOB1hNkAtXOoPVCS7lC+/PgujYdKUBPpDdusdgKvn8p2YJUTD45jT8ekzvsRAd93NZrrAwASY
JgRjSUdsBbvlFkBxv7fGXd1Z1O9ooZTIio972tfuZWbw/Op4TwYLvgzF3JEZFgXccQ+dmZTO4rj9
oPC7gJngExE3CL5i2K7u4FDRUUjAsGcTc26JFEDmJrGkegpfYb4KI802gAvHHB4FS1VdJv0CQBCy
Ax4jQJLQRwrtZI/uYObs8MYgOnHHT6C0YnjmgQ+7zbDHYrzC2O4CGQZRhY68MQCwqQT74tQSqCAp
oJrlO19lo2x93GWCt3Sps4k4Adq56Nh0VqOtaS+l9vB+r4j8G89t56qDd5E+ZXwkbrKLSlhD/XaH
w0JeTMhpzT7Q7U3sgMtDDEATZ5cSvYX7eYYtrPpw2SEd19FPoSLWC/lDMBhXJF0I2iWO3LljxsEV
wss9AgoT/9UHHlr/QalFOd/zSw/OYox9ON2zP5Q3RYaDP0btluHpK4lvpVDmXuOjTH0tn0DpRf03
M7KToU02YZVSeVV5iKQbNkDo6UfdTC1x7vrq3KeBShpzz+ehCzBtUyTbLtegAJrf+tpy6lHlabo8
7gYNtm/b2XOqsSRPTmugSXy3fjQUp2mMPFV7HlxFD65px8XbtIeSbNdTOFbi2XeWJFbnvxMCckiv
piy6Zo1e8EYRb34+h7Roi8RglMYy/yLX/YnvygAME4ZHISqU/qvlxuH6Z9ANZpUH5aqgVYIHdf/4
qjd2z1dUxBW0MiLk+3MD6pDWVtO0n8Y0m8fJjA0dCqSU1sPwGZAKS6wUhB5u3GFbEBaVLWAJ9soi
vjSP3WCnfNkOlWctrhs3jFmUU9uT+kIT/d+EsI54y13cRkkV9LEJauSeOEPxMQc42cM8iTn+UZfq
TAIYf6h29kGXw1eDghYl8fmki10q1UkLk9Zg4JCqI/j/68i6iyrNxjCteagNca0IPwHMPdr9QuyW
siTudU3JHbfuR28nj8K9+FhKBYoAqZz1GTvQsagnYmu6IQeVM9yMMRViiEd+q0u+IBnS701UdOA3
GjqAYcbVBqh4vfq4QfUzhVkwnUosrUJXNNHysG6KsicyLAIKjmastXKIKFc3hm1Ny/Nw/MfRt2b1
HpwSTFW4T32WTPtp2rCF2hsx3sCYTnIB8N1/8d5GVJnxXu8rC+G2ZyhFtGLxAG4UGJflZn/2uM52
OTqo3jr/ZcjqLsA08C5CBXSmhr+Ht2fOWiq9FWkQ9S82y1OBPrMzaLfNfqKzGXX8wpjQ8lYYUvN9
/pasydg18RYpwUcoPkGbEvqY5gPS8wURkHzM/0KGJUvziGc2qwcEYXqpYCBnS1n3QkmTYapVBHtl
AMqwy4jmBQN7BYOTpq9ZRL/qz3QHohYZN9+l96c9kna7qg4HT0baVqJDgfUtjNGSVUOJHvdtI6Im
o+jfbG15tIwaej3gu4IVLiJ3WNFm4Q5+defDLhO5TvrxBBFx+z/V343U3t1ZLqRtKejSEalYjfVu
efeT1nJX79fP45gS1jdQG+w2KIRwxe0XpZNDnX6zZxgrBFqEPWqCLnFnXnN2iKIPjxrSvYit+cD5
wwf0jDYpG8EyBJMZPCKVq2NTghC3ux9rOimD6n2Ln3IbGNBfwmxZXV2DLePscURJjB0cQ2qcoQbb
8F3K2of77FeVBzSGJwwCX9QQdsAFHjfAaa6t537qgZkTNIDU40aqYTpJF0WIi/AfmK43cgBtFje4
aKlThWCNy9qY4wLSUyXHtqbPkjCucZcBZSq6otADfBIq3EWQ8tqCcQKDd2fYcHyVgpYg+YYfP/Vv
EVPF4cRDgW3/rlpHxD/okpLiCBxIjMjS/hkMODIO53JcthAnrjs7/kM0KTN7wHTWJFIpUtW2S4J2
Sska56DNmcRnlywjX2s6FCE6syGRpUAEvpO2B4yk6VU2+XN80/g6gX2TegmvraZRXMR7xWHYJpqc
lCyvRXRJl+V1ZriZ9FYQCg+LKg9uk9lSp00lY0jwuBXA3NGXw/SSPCuRcf3tRELZui+WBH1dvaHD
WinTXxFiAN4xOEjiThFwT3f62PwFLdY7BgrA9zs4xf+VvJ7fyKZe3AfWAhtZfL3H9h8dX37p6at3
ALiP0/lNcJK+WWvTfvQuNxfBjCdLb5d2MT/qejP4mVBTd9TFrXzioAjMOuNY5TfhI0Jo4KpwBrA3
2swCM36/sLY5PoiS7uWIW9P1kX9dRUlSDURAJqOdoU/MtDafIGFltCArmZk3yxcNJVgcA5uGMHnR
KygpeA8NYDliRZlifaI8PLcX8d14h3gunpYpggrJj9R6rbgohtT/f9Xq4BLJayMbuJv4el61DxH5
Pb3TsPfVzaaIC3eiSwxe8t8B8c87qyJbFzWSvcKIsb0JlZ4uLgeyvNnIgCqL3xQNouYU7Ho3OmtE
TIawET0OTK9p2HfSSV5agm00in/8ID9wv3TtigxZOKEz3T91k5JVITVu4yzqAle/TqlB3B0qZ9A7
antuhHsmyn6mJnsyxxLEe18u7quYgLmBYnb70pPb2ts/+B/Oe9zSaWx8zwz3YrEPTQpuYKNIlv7o
XWD3QCU91llnG2EljTMm/67frTZtHkYk96Z4Meo6Kz3ONi9OYuPXYWiof01xrZy+JavxOTLPVMYu
omvsv2/ajdMIRHwhRvxVoYaFRREBvq1xZg3auazVaihLjx6dHiJZqYMLOhV18vOoa/vIYa81S+7n
5yiX7PJdwubsx8e1Jw00Jx0TU3gOxnBALhCSRR/0kDMGQg+w2CPuRU8XO0z0MBpLktOfeBymDSA/
nBP00hV68XyfOvECyZBW63bNNoJua77mojKmkHQqSo48XJ/WFrjwY9D9fempnPQCfUiHbJ7W69PG
waJG/KxeBfBJbl5hzg+2UriShoEilf3A08EhkEsyRDnADenlb2eATR1QZ5l+zcCPeCzRawyNLBFS
S5LkFK3mHLZa2pMHZFHW8sv5foB/VW9FF/p8vbvkaejtDiLrxS8EDgP9CAAHNCjfnXkDELLkWcgs
cRwbZYBkUWbxKqQjVmp9BWcfMLNEplMa/V1MP/mh+Xgfd9quH+VNQWLOyIQPkjGlxBfhA+zg7yHF
oqNZvScsDC4etH6YE5s1fLiOeEjxIeMZOIwQsOtrkOm3vhoStCvzVwJYHL/j1sg9aozaesJktD4u
PwzD/0brCic5016CKacmVh8kASjjL520cn+MN7EcqV9PrCS8s3MqxHuvaa9n3DyFNtbxcBvN/GBG
aikSoO0isCw9kr2qt8XsA0OSAj019XpopuxRUpYVLDu23WR7tNRXEhLMrxYxv2Lsj2hOlcHAP8QL
LDnz6H73FdvyLPO6ntjhqkEtA4D/AXC08OjlkLCG60YgFHsUyUF6s5iCVmqWk/nuW66jUoh3zTnT
3NC8ZLWQAmmN3oCpT19UOA0ZwkXQETE5azX7KrzLLIr5jHMXMDWeHEQUYrg2jaAdMuMiqviTVpzW
91IA5/Eq2uOV5ms1w2KPa44hlRNe9J5Z0SW/Cr2+2jNUxTxSL5abVCnaj3/1RmCskfVd1kKvAX2F
H+FD8a2sng0G+PjS08bnSXnlusY3XQd6a7y1IQwl2cg5S38jpiaDGBhd+J25Y0lhtRSLtRkAESng
FyV0ggjBgeVr57FkE3HFyeK0uGH8/inQ0tU2v5QsZl59rndaDAVoIIWfQmJHmbw0kybMNu9ERzIl
XiIQo7EIbBqFcdqFG35bCkjm6yna2vQQFoD9DzEQOb8+idGJX6UOL1bSrv19OxF5epPzXJK4yWzQ
34EYLuuNMJl0HWqSn1AAoPRag5JbogAVJGDBXwWFoIfeE8Bt5D5sneRCpmmppQI/BNG32LH2SEEc
6YyuOPmm8UQk+J17pSj6oP/OEDzrtY+gADHPQWRBbZlsUFxxJZ2ntjIy1TFsdcQs4gTXyhnq8Vw3
G8oDIDDCpF5yG4l+RSJUHVjb3Z8278NvpKKP2TRq6NFtgFpuyck3IyYvtgcAt3YoRk0aOt5R94J9
N7pmqAUEK6lUFDYk9V7CI4A9UeokCDZHKxt4ggWj+oQdMs0wayB2eKyBeP+PpXRlrr3NTu3MgFAA
hX+oWWFdQGzYaWi0+acNYNTulZ7eY4sN9QnUl45nsBCm7xzWpxLa3GA2hm9VZFhdjcKTiuUGoFme
uYtPGseZVb2rU8uORRwivwgHpWaZNJ20hkUMYirUsJ1YUpIdnURw9ETwshOTPCbJZWLLEVV+evA2
uIMOe73UbyQCM0rL5Qpuz/J5risHjjYeYLvAd9m5jzzT0SZJqbCDlWEJ39XIKp3IP011Yg0rq2ou
Lyte4mQCvhK2E2TCgTGrjiURai4h9a2MdZQjwrRaJn6gOX29lYLr3V/JN+TQjFyDigASlitRUpCJ
71JGYG3k9USHPndUDhXNfISprzDSG3TlvX/A2fb6osxADBWFlYuIXuFpKSp0WlgD8/JGvml8C/gz
vn/5XSFanE3CBE8eCSe0uuh8Bn08TClRy4fmrPyB6Pf30pW5j6bF3iFcrH54MiACrNN5sjYufpY+
dHbr9AV5xfXSB9dHm0S/8j0lUy6G4dn/nq7d/NkZ/+DzpRuHgdfjG0LwJXBAn00/6iXeGLG91obP
aoLUDMzaX4yJ8wwPpNPLOabaJM7+K3AqacF5FLwzJ+ucbOI4dgUXIB4Ajavggmuel8Q+aIxxHvOO
el8bfId0K3AS/uA7rJ86CngQGLa8+5xVNOcZkhwP4xKWjQ3nLr3k2CQHE2NbicgR3oYYytVOlJ07
nAz5f9abJBgN1gzLlhgfXltExNFSTEfexw1J593y2DUWHMBNbXbWwMaXY5vqaA9/Exjd2kO2REpn
SEyv8lYwiWzuEi0AQC/TzThn7gm43mdZp9HU/E+VXtXe+bxXOR73GgaSV/K7IGZeW18s7b9edz/y
M5OLec7ofDgREK/HVyFCHG7RCjzErtmnYbcEqDRQ4JwIbqo/DSH6GM7QePTPW38C1EsV+iWWxdTY
MKOP21njFY71QuIOCLD0jH8l8wiagO+aRDTpKaj97ggAsSGq8iulmmCwjugSGIB9kRXuOyIphIGb
EmUE8lf1d6UHGKTkJWP7niMA8KuaQ9tmQUcFnI0He3fMenbe3pZGK4ECZK6A253gC4wxg0TM6Wfv
g5PE0Ffo/X6w7k6NPSzllLoNKa9SDsNjVz9Vq6BgZtOHGG2jwDViyoOtg0XYmAmLt9+L8aQSIbkw
yBV9S147QTt6eMzEQ/MK+HPLeNeDX4LY31YOhtHnSc0IV+5IEMj2oHy6qw/lcPWW1s382Jgl9SNc
/Rj9CIpRNYqrh9iaPVjKC0L2q130JA0lg+pjG0KVOESoSLUzfWXqSPy7tHejJApStQ/jKNK2k3I1
HsPikqqaM7LhygjfKIpT0iBANY8RdHP47cUEEs5JLdrW4o+tbgBsE5jaqZPzSwtGICxbp8cYpCC0
DD7sY0nvAgGyFikh1h/PbIJBY9qQ7o3Z/TWbyFASyYfTwRZaARhFrQmCzoxoNHiM+74J+1rda3vd
X9PP2sN3Q3nuXP1a13t02ema5x7jDd4yAloZomEgZLt6PyxOenjhy6+t3MuQIbkOgRHmYbFnFB2a
OX/cU/8NiC5LxhH91OZtKvpZolwCPbczE/7EOYj6kCdYluwc3EHH6tdHd7EUmqwFHVDb1zilHddq
iq7Y/8FaiYZqhMXuqm3HlNXZwkVebE7wowWYUVWrUMKdXl8kOtb1QYY3jc8Sju1m5zRdhjNByhqW
Ochuzh87RLElm5hu048KiMP/L5NhOQs1hwRiAhmU3idzA+W5THh8vkgHs1L2Kr5PdKZgtI4Wisv3
eYoYnngBC3SU/fWlShE1EfjBx1W3ot+OsmRWbF8w9vYzHdq+Jw7TMEVrMjzgwEcfiMitb4NviUma
gvZ98NIk10GreoSu08TSEG2bGdzksW/KH8uO6D9QAlhNomKyCSWxbSyvvH9atoFhAFh6FxWtm8N2
Z8se1bdqRYkXx9VvpuRbFjLsMNwPJxHi/qsJlFPxi+jGyiJoasKQlRq346F5mwd1h1sgfVa5O7qh
Y9JjAAKmpodTVvn3HvSPPNYBxHh9WlJ1MfsybP070dcEcpxcEN/s6R0rF4AazOkULlMnB9QwB1QW
37dNtICvovzX/XpcpZ1EPHS/uInW9BVspc9WdbPsbmIlWBrQYNB2PVTOuL0buK3TP3KCVDw+1i0x
00vi++VmRpMUjd+2ozCU1WLgqEadgJ6IRsCiOhRq9lPMtSOg0mAiM3KUqhHB+zleDOgg11Ho+w0K
xt7VoyAajIUxVRMpL0wGxsFjDTwTjQ2S/24SIk659LbycvJt1TihQu6X0vRBUcBi0nJ0hPuv3yj2
PbkzEG26vDAdljIUTahLdOM8bkjLT3EF8mcVr4dZiagIRTAR1jIdxD50KnulfPpPE2oe1Jac3COo
7SVVerqhg72SKIvfFDsj42hNJ1FbWke16C7JdGNn2JhH02abTzD3H94hzWkVrz51yHbywadaC9mp
RCq4umHWRu3vgYNw53k6Sg/YwkQt4qEpHI741YqRV/b97KuxfM80ucWQbAFounotVKl4/RI+8Sqq
ebIMOmzRv174TDqUDnNgDL4A98CUhJ41LseWL2nOeBV55uChsjjkyO3lx//vjob8GddPUx8TYlk7
wap+GrRPucXDJ5XsEB3giqavaPgVRRM1S004R8tGOsetm79B2Op0XVjoUWFpqcBespiUnWCKKyMk
KcQib2ukyV7AiRIM8vnnnZSfG6bgZzRmgUxFi9AKdhvSlcUDqqFE09/HTW1kxphZjtUNmWO6Wg1F
5ZxJzdgHTXdG81SPJK//4wo4YYWivOn3/C6K1QeMq/Ip4c7pW/K2+sekdu6d70Du4feNEHB9Y8wK
Sfqu7cMDS7OryCbBLtJrJzQSaX8zrq6f8EyydFbp2tEaSRqe29hourKRDbTVGB/T9lERl+UZafAf
UgU1STUUb7TX/KjwayCiE+QOBeo3mPn9jw9OxE/9u9hxo9X4r7fjqiBcmJr0xuBHxaiE3gyqBim/
+1jXRa8jNgzuXvdpGgBBzuPvh7dtjefypD0z+Qwy8XhIizbZf9RQ+Y2Xfm7ZeQMkq9G9Rb72B0fg
WF/G9+Kl9ZU27AzKs6fuwsNmnpgrT7W3+wwjfEebbKWKTb1e2j9IosQEROUe9rMBj6nqGEFoWbA5
d1JLGCx1paa7wCYgzov5E++OZgRtFxRpEqxLzplSIoaoDPne0I8GvUd9+Ep6Foj2RukhefYpYmPP
tzMtptbTcTPyRLJj8C8KhLmiQznLGq9ufLrpnWISY66p7A9diJUuS7flWn5neeDaBzLxEaaSfk/G
B3cpcQwhDOjVDrCpQYxQ0mfBK+fBPPgWmtZ+HfjAZy9s4NUwnGE0e36aZFNaBoMw99ZQPRUxwmJg
yft91sqbp3JO775qCFulFhvPSwuxEL5BaQAZOeFk9Fcswy9yQrxgm279Q9CaRZWs+ZS7F7dU1nwk
jc+OYx+bpMmYr7DeDZjeUDpqHQB/RGTOV3ky/AXNPCzicxDgyG/r9x+XMDP1ss5D/0cHkPH9PEck
nOzs1EPGTZP9x8r6h+3xBG2bIVLKsBj1krPIMp4pxbGQS/eGl4e8wEBaZyGcCZy4vp5zJ9tdF4of
kuSwKxfw/c9Nrv0cCs2hXk3u7bF/3sO3EnuZJ7O1Y6NXi1svgFTgvsnx7ewg8l0ZM1BSeU65DB5d
i5y614jfOGMqfGrMcSraB1ZPk07K7F8x2VrxzPMW9bEf5tLjVaEOi2oPgmRzihGAiG8ybhIve7Jm
wBZbsfVBlECebdCyJ5ntaE6KRFDw1oVBxm5n7R6/+o8o2Zs0eRRjXvpMuux3g5GyQfNsU2vBCSs1
kffdB/1yLucqm9l5U7a2LfD6GAZ2U1bjuIzUZlBJo0JM4WzBs+rXq59DdLoLqdurxqi6WRFqUtGZ
VEB4xpz0BiX3nwlLVh3pXV64Q7GU0mrFVOSlB7W8RBMg/3US0G9XfShgClIgtXsmLGfQoSHGxGWm
EsoKBXldKrzR0KID0FMBzu9ZOXS2DGggue46tgien6uJn7CFC99/7OduiGyyp/WASUafGYvABrv5
H/lwkW81ZtBaH579hvLRQDDft9zTKnDXHvQVuw2qYRxTeKlVWBY4U7HiMm/N/vOeoOeTzJzZwdhV
VgmY6vO0+xIHmgAjpU5bazjCw7xlWy5+X4gXASD1B4Pikf9cU3pRqFPTQPRuhF8G6K5XRbalXCVz
2hVOq1OGymYUznTYz+JgZHgDiJ4OqHltfJK8QctBj1KZf39j3AHhN1JBGQYZluAVyOz8ss7bccwe
NVAXGz6k3z0RDfOERIEFj58crzrI1CpjIpPhsrENniL18tUeLHY1R8Pw3mSmM4Azjc/scRzYaqLA
DeQWD/f2mqkuL8FdjO51SY0aatZNMtUaLgI9TJ7Z4AWDNOqOlGem21h+teCC3B99BNApkoufx1ca
2ndD8iyafuqu+1b4xosaJvHDie4GuN6+4EFpYUXkPtEivpFtfpZx7P86t3NMRcAJox5S0llwRYTt
1mYJZaumuPYBKBgya0mSnxpnJJLEh3Ua8iS9n6vGZsndwY4u6w456Wo2FyCn2kdl26Sbrcm/bY/1
A1GO909GqkfVO/FbAF+V/OeJ7kzEK9D+TdEZS12aulq47fjKNyim2FoUFU9CSPCmydaXUQ8WqpVq
8yEFAW1rnyqv2wZaVRHxqKINUY9I7/oSZoidpAbWm1xTAIbKAD+/ccqWo2D2001lxSAHFW2eHC/R
fQTWH7o9LmqfS1u02mqCkp2alEf1hzkWbJm7gzx80I2FGAnQ5VAiwBUAl2Y3+TmzQxPwEjINngXG
Ir1BkSE8sf56iXXYWEDG2EGxg4gHLQoIr6Vwgtom/nL7n38B1QECo2xYsU4cy2osg2Ls7eMOZQ/s
5EsyDoqx66zIJ3Z7iNZ1Wbr12Zbf7MUtLYsI7qzq+/UDQkCHoMFwcA26NVRKqSDa3OH+b0BBo/Xc
koB8HnZ/YZDh1kJLzDALiIzzn5P9JeynzVuZVmzPdfAF1eu0dHRi7hDvcc1Pl014cxwPsIxyQqw9
gxDd72OvqWL20pTEjq4RHULfd45K/sWP6ZNKPpSdXPwMXNrjaBeTXjh/r7Llb+r268Ag99MgQQ8p
bQKYH9RK/4EJiyC8Cp+lCRg7IMBTi6YzV8MAhkKrCT6AcDNlGdQFHWXNR9bNlF9Mx5OzCfYi35tG
pueWa9SEC0ff6/tIFZrk6LpJ0kolhzxOOvqMNe4yaGRybVVmXUjvpQJPlMIPg/9fITDARlP3ujSi
BrWZbhBytr/JZS42VAv/Slx2R6BfnhJr8s3cq7D44LTTGACgwK1tjmAOY+/P6wKevP7BWUb6aOz1
FXHyb1TfvQiAu/YNfk5Xke8sVHhzr7fz4dxXdcUqpRsu1BynEz+i2xcpEfRnC8Pn3yu9iC1AGc41
Y9iP9l5ypeNmkhrVcx+I+QLVp68/jVM3KSZuWJqUSxxKUUv05Fb3ymHj7SUldcsImVMdxlyJgBAg
PeY81Vm0+Ar5s6/sAlZt91GedCmyMQrQkIC77C8mnolznvqI8r91uMz51peN4B58jzUE5AqjHYAT
GjIR4rIZFZQkvD9SKjUXImoyBRlVrVNCM6Oq6WZhSd3WECMnkWFPBoQPasvfFaJA6qMdFDpnED0k
2EMdSDXqbDpZlv1Irxv4G/BaP1Uv2p5M83rIXUyIWTg4Vcc8g33pvMoJCcnghXsDJcA2vGGF2a/5
7nD1L3t8l8b446CbfYtSQr1/K9SrBRwsPoFG1DQM9VMgo9q2ZwFaxnoXznFAfeHBR6LFyY9oCyjd
151F0pNu04FBBekreVTpmsMtnXq/gAv4cQNpdxgZWhL2M0jFZWfrlsp+QBQTvCN/Q4WJiQEnvHrW
2XXwqvWX2JXfBJ71YHHpaUfWM4lXoeaTFkT3VhjK7Zgi6joChWuHeJWkCVbXpzmwJj7TVF8x3tCr
pIEBj/pNxIu0T5ILe5YahireYbhrZH17t+lSrY3dVeajq0/I5jOfajc5gPCXjLJWTNh/1lZVmUt+
S163U5DL0FFcmQKUV9PUwPudztVTsfZC1QZFF1zFiNfRiztSLiOcoRhgH9JIRMH60roxmS39rhJA
/zz5MpqmqFjSlJsL8pOY/5H2soisIJtWREk8gT69NEyB940S1M1dEgbW+VLkjbOL49ekkTo2Yat2
RGlxyKvVWwAFrGNc5JxX4KAuKv0NYPjXnYqkTRwNqPFNLeaYXlDn36kbMytvb625dcKYZf8a9+MG
5ecKtBaWoSpEj62lCR/Qn8vkRiOTlCI4fssNeia0LPS52ocUS9V/EkwSAIIsjoZb8ZrcWN77MKsH
ffUrF5/wo8omymfY5c2B0p1Ulppn3K1fhGdBEfEk9T8GEydWD6iTXBxWAen9DlvA8ofk/2rGK2Q6
hXRbRv1IVkAWr2iJU3NkTaBlecw575LVJBI1kRb8CxgeSbOfzySlIuoZjt5yYMCQ9xNpeRKVg3q0
lOsvqXKHTLc+J0OhdGlvef7KlPjwf+e5xFGuZESuqwNUxjXtPvH2Uqe5Qe52nb/rrKGlf6no2LbB
C3SK+pmC9vsBOv+SaRs7+J92dy7eJzKnfAX3zAnxk6Rt5BIFrzlFKg5UaELbFu+C4tq3QToxv+eU
JID1A/zL/DKK1Y/GS5j4brvMV/Uf1ZfAUcehvAl80N9ydwqO8EKtAAzlEEkSW+iBtxpT0EooI/Uf
W76tP6m3eKjGBd3kkBfs8PNkyZ8X7f0a1IIbtsBsTZbuE4u6tUMJuSXojRXgpp7zt+lSsa9JJocN
YVrIXem0IgMpEaj16sVaZ9coBbPH/ZAWH4UVhnoLklCjZj2fAD3z/MmulzusXEMMOVkAsi/LSgxS
pWt2B/K0kclqvLK3ai05hw0tq/i9rq+sXFUmIyM+kqxCd1cBKJHsYuCtBmPKRjMrwWeII9tnmdOB
bmXmo1Fcz8pxZ/OMCEynSm67HbYXlaur5f+hncz8zXWN0DmBGZBmBwqhoFDrSsZRjUcfY9kCVfWt
SwP8aFbf0TmXj4uDMXfERaAehQwLljLk8CdbXElJRPeUWe8laz2ofN9mkK83xUhycD3md7wAq0bl
9dvJgmhGvownKmVF2t4tmN9wdH3S0tI7/1sc+8TJHy4JD/O+M7Q6JAKbCvH27S081uV5XjmWKS5p
AzJxec1e7gIQXRiiyF21u5Yl5EK5ueTT3W6rTckL1rJw0EV+1H383Z5cm2ZqbJ6dHsqzjb2ZX1PF
OewdjWmku3/xiG1qdw2d3474xqz14Ml3SE4T4cscrOjCMjV1kqnzMk+//ibKzuUsHhbkCcvfTOKe
oYvjXEHAUW1Ctpwgd6i12NdOy1tRQH/BxwNyq4P6S9sz9lf6UEk0Hz5cVpPnUrloyl91y+0bTWYQ
jMhM2lOGThTDLrVQ6jmR9pf718RDMVXGWSsyDn5KSKgpOGPRZCO1Yd/qKL1yGLZSXbG9/CfrfW1p
3yqlBxcBuJmxLlp56QwUNKrOckLNbm4dfaz+VF9JbZhzIn8/DmfG+7xy7AdXvwzFc7l1IKsHF8F3
FaR9XDwdQzso+spvRLWbqf36wAeiRndNj5jMnH4uXWvm8E9CCCnViHyqgz/8x921sr6FNCYNNxaj
8pWHZDlN2XZf7lRBpPMLjp1t4wJ4k4PnxIG26Zeg/Nqbf0vw/hnEu8wLZbGDYfc719+/uOIwd8Ps
2AbL4WyHfY5tHOSJPMDTDNUqcoFl9VGY7pO7KJYFzXQh21LiCvq8hsLTm/QO+NoDflwCoDYCDguv
bYMrUf+oiVo0emIH81uHrxzB8c5ew+XX9Qdti+aoIudarpZxgODlvg0Zv60rbKaKXa0M0mB0T98J
YhCEtzbBi0kjX/q0eMVMKy4lb+1uKMtYy6kTQiDB2UX14ZtmXCEC2kJDQL30PozsEbLGVB9v02Wr
HRgrRSKPIGfgfZW5icPGUC8v2v0pB2QxuGt2jtpjy5FAqw+VQVPRCV8bFimNNNX+/x7iyO+l+7uh
q3W7QwkDHIrh4UUVwu92nhMfs8boQU9o7YXMVM+aO2ewBI84Sh/O7zVCR9qSAtVFyqxvm06QmvC9
O3PCVl8fKCtHf53dXlJtwfvAPJB7QhXQrlS0rpHFPPZgeuUGwvseE0wSQ3dAxWED+glyqNVi2CZT
31aR836TqlmkYr5g2LLNvsk9AXgru+Ss+2KUoEKYTKzgLAFXprn6o5O2pmPtjHuzUs0uIm3EFjJq
LrjpAhuH2cMpFM48s47u8KtT9GVS/q5lZct/JZ7scvUFxK7acFPVJV4/+ULEb2SL67XYO2mKc6i+
BEg7TJmKB384MuAMxe75KSmBy7z3H86JybVQxtZwhCs4l8vKmy/pXfKIos0LCU0UXp2/FWy/+uHn
pYxIHkzUHriICBllL94x7MTVUb0vc4qnlyteCsPp/aC/mmHvAeX9syTAiuOYi0ViGEFgb8J6nLEq
NtR2zcxE56UmMzlHrQpMQphJVcD6O4F/856b5ToSKIjAqHXD31Y+BXRpJwmzpNFr7nQSk0coMBvS
YjQ86TC4fbeyRM0t/ASUq0mG4BQa8elgu2/6GtGUPaneceLnHBzm1kr/TIO+5/2tCt/StbVFf1Bn
JqJ54DLknb6ackHfL07ThyA8lTlUf2WtoJZ7p9IKjWwXkxpEruoRBuSG0GEMeINXGo4NK64hg6e8
Jv60q/doeVSiM6tCEN7c0tfynoPWlBMbtKW2PWnsqyb1DN+ie0OfHW8TACuVra4H8WgNAjOb3DFS
KShJ/SwM6jqGkStIZV0QI0a92gJy7yxshy34+9p2oskT4yvAulrPjlqhw+FJxMd2KpOZMlLxKVCh
aS4kx123OzDP9osRMw/Ev/DQVbYvDkoagewQajdkLKfDeHQRuqBvoPE8G+TNz3Qf1PGd+bqM1oqt
NBCui50kHC6YiKDVAtp1aaeBh8utUIrj16PHkW0Olq9/3fxFddGzMc1nwfwZlfx5xm5Fkf3RMbYs
0qjyEFJG4CnkMR66p8LVCq+5ylTCwmo1pAXHhqhwRtA+D9lLkRADWwLADZegeUxZWrDoKaVYR5sJ
b05EYw2oKwY4vS6a6ssscvUCqLJXaipKqMHzXwWbvpNvqLFz4RFXImJyiT/ETLSploYT0wOn+Wct
Z/cK/HMMam9i0kSQO++w4Fo7QtBlp80USorr5P3696eFDZNWoiybcqdSIO08mDAN7alQqJv6DxMv
azD/rsQTV+9QoRHg6jWjY0VOBaZyFMpu/XY11WUBOJCTRzovaL1xkJyRwPbq6AoS+jXmwZXGHFnK
30vCQf+KTokbVFllFPoDGvvc5lUhUgJUS4DeDG4a9AaPtuszyuuhJZ6BQD7YkKXieUI96G9M1uRk
FNX6V+sH5t1wehs0ayx997rHvm/D6cWydkDsKjZSi83EnNFMbKmJg99tkLmWhjRtjhIKkCzmPB0X
PBipR9OwWcCxpLRaV+9jIPSwmKNElolGWtAHQoT745fU4OwlRv7nzwDl7C4DdsYXt7RVIhamlvIx
hJJhA2mTsLOlFl6nkDPfJeScmG4Ar45+C5YtmTC1nYHr4NfFDbnfMIxcGZG4BaswVeQ+ez5wiAFn
1VLoh0QWaiHstHN4cbED1rPFvREdtNebiXSZtwXwMmtSTjkRX82pqQ5H9UjD+QWSVwUIJEIuEBjk
Ou53HppuP4J/IUdnYsC2XU1CYYSjVr0Ha2P+buYRMjfWlJ7FUlvR6eMtg90RmpLq+dkWuwMSQ5LE
uqbLdYbp/cklOPtndsLjN6eN93h0nWNCsmovXg2iyyvij34ndvj0JUDCbn9XzT6BBn0USVn2T2Ny
F8g6vtybEqE4shegHvp05sHHvUF6ZcUSTKX02BRh7A1Q13lV/c0BIY0iJPpSP+OY1OiqxquPUaGk
/v4c0Uzc5azo5riRa+p5oGM9zWx9IjhQHETjNIoAGOhgo0a7wETZ20bfiQhqEqdQW86ieefQNGkQ
MmPJamgxbhbPm7mPAV23iQ79o63BZsKnnPuHlPu/5Iw7sX1nb3qJsVSVD8Q4JStMUzb0L1ns21/N
JIK9wFq8O613hHep52P21Di9vS7NhaM2yu7+/zIUEtr5JZkM5Fn4I33lXdAHK1MsasBYfgTvqx+R
zCMQA1tY8gEKLEMFBdx4OcGSvS+8FinltiFHL++8XP/ahPQP8tiDJni6yycKMOCobocA94yYYhJa
dPjWLGwgunxBsaFuZLLrt8hQAeLkNhjXN4eQN6rtkTX2LNdY21t3sdol/M3kw4ymrOxYKGehUvZp
OUZQXnyt4UOOraG4EP0Fj6EuorD5qwLMqlogyvZOzta1CfPlDrJkVUQUDgwVnG3ZBi242O5XshSV
JPyCu1ybp8CO4ME+5QSZubyLAI4WXvcK4CoGQ5R1m0yJqoAc0swuxC3KNV/dMn/qrJg+v/XmSj8w
4lzyKnv9/KD3X4bKDSu9t/HiG3qeUKabDT7a4uaBTyDQwt6G7G3gxoUYpYzmkgezq1TfaEKUJ8sD
rWRVdK9JhHdXL6l8d36rO3UBwDqvQwyISyq7ZVyXXNGDpKaXJC/W5T1dEb3ZFAMrlHGX7temaETK
z11FUjb1ykfg5L7i5kXvGGhdLIk1SWj6gfCgtcqFGh/7AoM7IiDgFEZEmb6H+M/jCHoHCtJ9Xxut
4QddG+aJt1wp/5ah0mKwtBleNXXL5VxJ3en+kn1AbsKo/Zf3OVv017LDFQy1ip2t+tvvarP8lemM
HBxUgUEXPfXj0qwp6BWUG4U9762PsJCAq0lRfwbWD4Vl2ak9o6J31iQJsLOufeoymz/3T1rbrWyH
0Lywx+IZgyGhmWr0FBI3K+jTtTmzOPNsrg/xHmFFGv0pbe42i95tPXCLKiscisKL+6vRub40v29e
vgLLGxt45aw7n/5vPbvgRopoTLXhkRkzZFDTI/EADpjT9R8r8zgHVyiY+oMOr5YRb0SjaVw9gQSA
xbLEnJjD620x7XzVKp6rxIx+PhxSTWQRQPJYn2wiYE/HiqsBfj9p4vNuivrSZxsfqCMJlvWUeNqi
gHpx6pFvLixkVMWDTbuLKIjhqoBUP66CmEtaiQWrZXstdgTtbmSRBAOdp1wdrk9OGN/qb0zVmh/n
wzOQo45gYIq9afnm/0JRDR3DMqygXfuBnXdKAQ4SFksySqgwV9C1Z80IOwvadMN42su92tAQadpI
rn0stzt4PB3iooaGkqkcaPwh6Wmb2HYhl9S+zb8L0Xg3984n7FdbZKJfhb1OMFnvjClUQ2YCWL20
cMO5WHsJqbLOP1v7Lu5xHXJ75xMGU2Vt6U864jHyfgGRQ/0WaNnyKstmC35Yui9Kf7q5SbcHfXam
dQ/bjsM7OYf13Tjb/slllv/biKsqw51zEyU7+MYc/EBZY2LaTBu2BOlYMZ7eH5kqgAzd+Upl0Oo/
Z0cVZbIiQI9mqpm8eKTz45/q15kWQDj8vFCtnSrXATUIs/UPuMphF16NaDH2kx924gZ9LOWuCU4d
sxQ7EeA2GaAVzPHjcosy2jAltjuc5s1gy6vaAWVApLpCbZ9ofCgDT0niQeonzj3vQ3yyhiDhqDns
spioogRG0fciDQ7Bj0bcznSEaQwrSDCZpUZKCKIfonFM08y1uSqSmypsxhpKdn7/9iBwzKKvpvtS
kyEOAtbVwl2w/xGojCtxk8BQFDTOYGxqKA3d4VJVQUfhlphtc7oMo8g9jnHguZqt/m0SJZ9Lc3lf
+SNtPG62Huo0Js30+8MSuHAN7JJQxjJt57gskUjeSJpm5rWm7K129CGPNrXZM7lDtZQrLUnS8Y7S
feSDdArrkKPqi6dK+N7bLE3xW900Ez7wunGHVuOiGtimAadTNTiRaRTOg5Y5hC02g+HaU/0us0jY
EhvGv7eR4dP1YHxl2dSGRGp7D4qJeBdAgIKBssgvxmVHLFYNmwOOf1txuYjt5XfZSe0l2pcPAfpS
BsPTVjX/ixuNFQi+UjxVGseb2SYrzc6OHrGg2MMoXhqSEO4P/IV1dUt5n0Q9q0UQX7rT7VBYVV+8
O813+hhcvMXtjpb+V0tOs3q6fUfiqP6KNioXK3hec3m7+MGSEpmmRze1xJvKAjffE5CpzqMZRp5T
7giwqHhCACsEX9vXfuFEqnvVgLeTtPCAPsI6mj7VOXh/vkAQcg17WEtD2O0m8bhXHKGzC2feQ2DV
so7RQ3TyD9zq+eD68b5gI9ed9ELZYmhlA25VGHM7g7cnCGMzR11Kn9dcD91ps4jNpXR7bZwP+6Cj
yeQ7qRF/EJo0+KTxPAsMXyywWVJSCCijoG7peKv6ukRHnf7ebZa01SWw0JCYqw7lkymREcccg+uO
/OJqX3VlK5SFRisyyfqMABAPeYUhmol0xQY4X5GOnIkzj7Ekxaq+/aysqwHadohJsRp0D25Pg/1F
b13FJbPDlKFQnv5+Qarifp1dWSvfQUQFciqreJLYwu5zbs1794wwIXbOrZl3P7jzpxkVgEX3sSUm
oFqlMJGmyerSh4mX+M5+/IRlnppfsUwSOj/DSuVE65ULj02n7+eyddBw4TOUahPQQ4VUZo0vcQun
sc9Y1hDX+6+5mUynjyK7UwO9mbdWTnXDB2q7lCw9wPPd31/7rubQsmf9sLdvvaBCbM9K0mmF5Cn9
cjSkvl7T7sOK5OjO1HiNCnVrEsjiHsZ7QtTUw4AQUVlBaAS+uKkdeNKh+D+eMlePiLEY3BFzxGS8
gd1vl5q/UETfCUFaosdELWh7imRb5rxhVRCo4+aHf3e/8w3bYyJ9KECvCleUCTu/IRP+5wLSf/kb
Pa9w0U6An1PMldCpHakbURko4FW4np6OuriTdpT5vQ3cRiRf260xu6kNzGBKNf5IA44QpNYuoo2b
yhhXcFMpW4p3HHiOvYjVU9AoZnIO0RuW440V1ZRRhFjTyZfUUI2kpeg6NMZIGzEKn508uynhEQlm
2PbeoC6iudvY3gC34c4TdgnSVoD8VEH/Fqw8/Htj1r5Fh3N5Avh7zXB1hbkXFuHIfwjW12MYqPB0
QSzS74Ve8qXOLyX2DzozID/OAYFfH5M0/bI9z1TkJyxojK8XtiFhvabUIXRXajkIvM0/xwkIgY3e
USBvGEnPLTU+PfXL9uZGty5OVEfUJ3oRptl6ruannfxSKK+iBREA/Bh9NHQOiRnL2lNfqMX0r6e4
V+1EsN3krzUQEAewwp7YQlgZdzXEh/x5q69GfsesvYxVy3w/rqnWeK4SgFHvf3XuFsbKkRqHwAMQ
9AMI14HPYrYWKNmSlrx4+5rqiR6suoGPDaVFZgfv7IkiUupnWNalYbv5kIBJTL+GeBSWbXFBDMAq
gtdlRtjStY4GbSb91U0/x1ndccqT5+YJ4TEAYXhwwyivxulsdkL+kv5OYs/wVps14RoyLzqL50Vt
Nwz9ufn3QNQNkXBqcJt4WiNeL5f/FJms1gFv2wHMJiti596y8MUnULhWAfFXiA4whKsUQpKuPrj1
qMGIIDmqmRs3fASgjHFpQrHKtzQnpn2TJXv+lGP0zRrEC8OSUSoulv/3QGSrQmufN0opG3ezeoIO
XuHnGJWhIL7idhF54Z40XIonYGgI/Qyf8dl20u2g/MzXovxB329OzkpTDJo3mOYG141ktbAR67Js
2hv8unU1QBqoNgCFsBiJ8OG+8e33HWPgB+Us8/4UqDV2rUY/sN2oxd60pbSIgoD3u1gh6GOutsXn
kRxUDfZ7t+35crxPCM0ws/2O/wN/djyWJESp46d1Ugg+94gkfFs1btDR/vTSkL/cLkVe6kXUk/qt
QPGlPtQ/TlB26R2BX6tWuwN3B4xK9way6UyBYSAfIfu+4Gq8FK/i+Oid430nN+cXEbkSza4TFl/7
mChOZPtHhvAlKa5xr7WXo/+Wg0DBWSwF18aRNLJkQ3im7MvH28ANPBNmXTrZLPG0uwEbJrA83Xhr
CuS60XuWI1/MTVyhjAKZ+JbwKZw8IyV6lYf/au3IojEnx/9FBWIhHO18rffhAxjNlCvjtgpeLyQt
bFp5dA26Wttaba7P1b3xc8/zkUjrRkYdbGUTa/LdVQChIKnB+0NpnNtb1/U745P/qoujesZ8WHHR
1oD3RAUFVEqpejojWi6r4g1nQsGTRPyuYPKy8CwNEAs9l5dBvH99tU82x2ib5nSo9u4jRnb3HLw8
4gkHvlttlRnoVBDXt5ntst3E+ozx6d+3VTWerRjpI9L/1GQLTyS3u7npnSluwmqXGmVDnbbZitDp
QWucx89I9wlnb8vMvlwuNnHE+xE7Ct9yOsutchoLCWHl3rf381HzryUgRR3vJN5sDX+5xONUHah2
bn/U0OB45goWufKYisaMcJCT1iq0O7hSfvw8WdhRlZYKcElIIl5zzJRRXpJt2YdJuMPyjNlI/Jq8
cB//jwu6NgAvYccTPGXE4baFtU3ur5xHGYCeZvmr0qdoO9vIg/Z074P25gtG5rTCs95bD+89TLQZ
Bg/Ub1sveAGH+GF55XGJ2zSQvFqUL5UDaGRgDPDzJ+hAR6ri7gxmp3CkukyU7VjWugWZcYFRo4Pz
2ewDc4uoytsbacY+Fw9KCDaqffb5lRe3kC2bjvdgNXllf9v2Th69LifUw3V5CYM58x7szbwzfsCS
j9CT0dgN7Bdz0t+Z9yY/ctW8oBChKueNOF/lV/J1bmFNnMbKqR9SxcdSK0+2D5696wCXAsvl/hwO
+7pCy8VipRhlvT4Io9ij/2042ddaNN1yW56GD17JBmVa6OvJuRYoSJ/lOXVOKhia+pk9y6vobqv9
biZ7E7g9r5MxvczA7qLpdKYXdw5d/07bWbNOXZwir9rMB2mKWTxP9Gl7ikQXKCjlL3a7qqHuhZih
xvw/cIGAlAnG4DiN1Owce+wSEesLDRYWLLZmztjEQ5KqsucxN2JtwUNXL25zv+9OBL/CPmxAUMG2
v1KeIteFMkjBaU8251DzQONyWhgdFT1J/TEASYpPgAx5Nyx/SB30XlSQhQGwpY3OsKWmhrZdsSQ4
yVAoSvVwXIark47DXFwbfCnpyADvt5tGo+X3KrCCi4ZaQ6UAlHCk2q8Y+2GCVlNQtao692pFrepC
etoRdIGRTwAz2X4XZXjGRJ2iUcGjPWbDOGr3A6thsBa1uLftsi26boBfkK0h6ojFoaK0MwmygNoO
dipvGROXmbHt3PRsACtTiXX2EWXKlDJx+XGhYRSqucJwAHnaNGV+fYiFpd7p4TAqTNLVaFli9wR1
ziQuw/upzZmaGN0DM5SomZ4cfhwjPzitgkMwdqBHNuGSX5nyAf27IxaB5849Da2ktDZC2emcVMwf
WHXmb8/dkJHEl2eRSnEZWd6ZvA5BNvxXsFMKyRfPBM79Ps66ol/9YPwRBtnyult1mIUGJTTDw0y4
4bn0ttG2euzceXwcXDqzHUVG9ZdJgHwOWhtPSano3TThIt1BfrFPAgjC/g4sOJXDCY6GpqX7Qsmk
PmeYAPr0pTM9Q3ut3maL0AvKNspr21ApVtJ/WdYAw+k34dJTYKSIH8lgFt3Fh7sFzfS4W7sEgCg8
ef1O9Bk2ZeHEeZEfcBMAdbRbJI0qyubDyQ1HppQYeSQSFXlRAYhM9wbf67AHEbArrQfP4ow6a1fb
bu9nnBjK8J7yA/jxthRVdxuAOHZnVOkVrvRfTug1pq7tu5tbxfz80krUzzkkAN94mdL9MDW97zD9
FlxCUWRn0e55OHbXavodT2zz3Keym7v5LK/tr3jwEgJxQB/J0R78vO3il53CZrjt1PLKvtUl3nQa
P7xD2p2nEAWd0qpfXX2z/ZZUoxWadYHiK5CA95Uo/POP1SS8OGgjFYD6xRZvr8sCoAy8083PBUh1
+t7B6/1D5ealFS748RF9Oawaw49UhGEils6RtUfQ9gSgxoM7RLNDneFeUbNcjbAKMpI+y7Edyi8L
DhXDf6Tb6SdaRiOGU/4zGDBG/f1gxOCQ+kcwCUbEc3xrH0q5wdbjyGmp2CrF5VYK3YKPAVKPA/Jr
to+REqxxjByHZafGGmT8QHelclWv6r3i3ig7T+2ccfmGzEOJ7yOo2c5Noq4J1j3+CKUuVkK0J2uK
SbcIHIBSi4WjuL6ja4XF+QJW1xp3Y7sXsau6bNH66qkk2L4+zhzxprhmbzxA3AwPM4uFfJPGTBSd
zRl6CCvPVX3iMhoAcqtyxj2ul5c5OL3RmNWhin2OzSoC8Df9TrFdzq6yj3M3v84LH01QeySOZPbO
l/+n7E9ASqHA2uD0iEXsNMfhZbW5BNrHa1bauj30ObqsBQuwM6tiZT2Jq2wgP8lxnXLHLyJiT7JI
BXtaOfTha9Dv31qPEc/Q696V0Gvpqsf3aYSaAlkK/yZ3O7Csd0njBY6tOdko1Hb4tnzPL5bAuGFO
A3k7HkH/c5pmj/HG9wwwhL/Vs6i2Z80KzaR5cbPnn0rnjVYBKVo/PxfzecUSyOkPYJmHfRJjXs22
WOhZ4NnI66S0Lgok2QI1MloMJN4x/F+pnqjDbvTIS8YOsX4FN1Q54JV1dfGCXbl9es7oZAVxe9Tn
uIPUu9kNHIFFlx7Bf1rpyqyehpHXKpZ9lGy8dHf0poPFt0ypNR8pvGrx50WC5FmEQaXTVsGTmjch
bJJtSKAHAedOcX0lXDd9vJ3t9pbziGRkx6zM4JP/q+4HkzcYsuOLlwbdzl2H4HwZ6yTGKpLStNiq
J+8fp+xAw15f355PqgJ5F5ag9T73SLF0WaMNWE14v/pOcfHi/FYIa/u9cXIKiPNFji4maCl46vyP
ggBrySnimCbw8NErts6FEZARvNR2YvxHW2nmC9i88BX7qdW/sGWMvV5cV4wxOtsKDIhepQifjNuQ
N9Z1FZ5zMaRIywbYHtr/DklmKnm76Fd1KHUyJBIg19OkmwnVUzs2JBEH1x0C9vXxqMDXUZgq8iG1
cd6PrL57gQo0eQJYAjmtGDLEejqP4gsQBbmSErl0wvrgNPMPh8L+3u5t6UHBGFJ4O7Y60+E0OJYk
wcu5fPRnW56h2B91nhBlh6x6M4sOzreDfnHF9MvcGQ5Fmi0MbG2R6Ls9NxkfZ9STDfI7rB2Jt9Z9
RRStKttYAI7vAKLxqtwU600jIFhQFXjEEgmUnRcmWSt++oKZdoZEUhp0wjA3k/IA0qiWOH38aLs0
6NG3KMZluwdSxzE8BFbN86D12bpBl4Jpm5jSl/1Yzq8RmrTiZ+z9K5cLey1M/xElr8rJGgUc83vK
rtRbtCT0+EHcAFi9XVTgPdxU929sBQ1SFbi7/7/pK9+8LN3WBMuf6jc0vIVtY6p1FFdMisXQxx7A
dUwtt1/vHrLP2u1umAVwTBWnuRMwkRsBWbd28GM4stDhas2ada2HqtUqG+roKhzQ2/xuyTMKJwKz
NT2MYIVqCe44/Z+ST/xv1k6CQrbGJsaoTP818XaRTxjbsQz2Iq/VtO+z0E18usFay6yQFOGySV/b
CvyR1yb1y9DYvo8JU7B5F3nFhEHikoJWZX9do3Ff2AqKGohgkimeYYN/ZrGzxFiXfv3RSKSNnu+0
e90a51aEleCEuHGqSVJG8HVQerY9+b/VjUQKzvMTLh7zcEUzlXbrAKcnz8tjPo/G2CAfOs0a75B6
QA4yOGz0Egg0GclG5rQ5KzCG8DPvGsvsumpmYHYXXdwpn3zvvEk4PN9SeT3CmQ/h4MJZHvm5tJhY
3njR2n7Dm4+20HQPvAUCAJBKJ/lhiPCCiujeU7lw9SUEZYuHqwGBCtwnhjkJKVMOewvZCo6iLLpf
axxMHXNau9Qnmx/cr501KAOb7Q/l23jrKJ+7BpOefxWkbOYHHWrzoZrHF552fG8RrWMVWaytHEn5
1f2gEN83dCpXRh39Ks8kuqJ8VAPv2GYT+TQaq2AGSlEf0QbRg3pO8TqRslMndOUMrMrsAauOYsTk
WHJYHA8e4SN/zMEc3yNi4TbGn+kqyOoLq9OT7RN1pIXhWvQrsQb7YMMXdXE4b215L4A8v2Y3hxn2
reRz1s9cMR2Zio2TuRKvMRLPUJ6IQfjegn/NR2Z4yO53qGqNV98QiZy8gezbF97/i32c57r+6XoA
yaWwpgYhtVz4FWZ9TxvFvxfqMSHYwV59hpDvNDP0B8kTizd91/SexbsM1eyQn+VxvvF1C95iqkQK
dTAzkBhNphZzmIXhBgNHMEboLAEmbWEY1/IEXlQG7VYT7hfE2dEDm0dOyXs++nTw95c503oymo60
gQwcM8TYJRXXdrcRrXhXQ8LZ8Acos/Mq+PR3V2YDRoNgngRkkzhEFvsUwccfYqAmubHASWsOwNgv
2PAIxHpDqapzE21FAjfe6Vh7JqEpNZtCKCwhGRhGOiHBXLRjAiSYmhIYPJgJKldoUvY3w7tVP4wv
MjGfi9KJmA4KyEXHge7kdjn3+VmgofdWWbFc3VfGws+R9w173ETnzPNCsD3BKGBPwPxJEJcX79HX
6w0e5yYD8rSkRiMmN/8RL6hk75Gqv/kFsYjRqlVPU3gCHN5vXMdE4I6OoZmC6Lx4OlkVVZyfnV9W
01Gf152+Yo4QDSvu6oGfAD90SHoSQ+LhAIam1QpuswitZIPFSn0egvxt5uLONl0jn5VI+orl+ZDK
DO1538TnIl0BokNbzRBeNxXFknAoEYVCrgtEAzTCahTFOpQRwZq+nUfEWvIbqyBpUXS1BKAdzjGi
NmU1wKGATctPULWj0YIEyjysSIeE98HcJoVgpfz81R7JPZ8xfYC3cGqfmjzmLKi6oZ7VyWJm9QeC
iLOS2SljSaeNyoOq2k0Ku9sNC9T2ux8oanDLVxSTfa5VMeXWlhCQ07IsEPz9JGzmOJWDpFd0Pu2l
Ca6Ofd7MEpxsAUjfisHdXwTT7RaX+JCYMqt5sscu7X+uwNCvvuHxEBbs6YnsiEHWLIXCb6K82h9m
OtQ4mmjayRjxwIh+8pHk9mdWGgStiSroDMd1KUwsh50h5CdSHULuc1vm6g3+eCLsAbArbzgHOvDX
AklkBczMRuWF4clbBe9rNPXCYiFjTif1ASjaQ9OcXiv+4yW50MsTeHDHMTjGiJqI1603+IIkzhpY
UEIpb6CB6qvTGB5x743/vPcIB3ZvW4HLD1RP4bzi3Zs3lyWq2N5NVJtjzDGavNNe+Wn9WuqG7+Zw
PS/g9kMioiLLOOtMgT0uu20GMF7tP982kH7SCR6V7CtU+xZKegvV+HQC/9kOuNbn2yNo3K9yprxW
OeS8c29uYXhpCsW17aUZQP51BK3j+t7gDh/flFtRVwzj7Kce/9uyd9XDqY/bvj/0YsC9D5bKUzK6
XQLGskh7Qz/Izjh2RvgTwcttLaYEMUwreJTeltKkuz6cKzGvDGvSQsvVtgI12AB1Jusym9ymMVOP
7jZKLIYkbMmdlXaDWIz38NobdBLtCSNPEUv0og7PqBVfHknaOjMJng7PmgW7uMzD1dArWcuG2pB+
v9ih1L5psXMzd+kJ4tcsgKLVvKwwjVlXjOUx5h5sc2yOY148Npc2waVd5oQ2LCgUUjGH3vjW9N0a
LVNRJfeGzqD8y7hmjOPGG34A58hBG5o/2iMg5qp4sSnGbiZxgTCsdlVnuja5J5+MJREguwDNBE3z
8jOdLHFvUpqzrbyEIvnS870aVbIZVPML/lkLVkrhVM/ncExEEt3YmhB9reZISYkxAnbC3Vui2zCX
qOgx/zLy+Dr1egDJ+8kjkxU5EtYyx2v9c8UqLZMgrwqQlSS6/Rd1yD9Q+zPo+NFLl3UvqhJ/soa0
xvesX1GnDRjJa+I5W7p6X0iXFbBvpOEolwIlc1vVLhQ3PgDm+jmMroYakJqNG5FJgu3A3ykZOdch
oB9o3shBJX0Dom9Hx2mhewT+JRlO3AqgTWkR16zgAB8AcfNEDWOQsgua4pH0V6X7yMl+G2b9dRER
XIEn5qyHVPYBHmRvw1iTKyH9V3QMyTrOa2nco+df912+rKCoRR5Z9AuT3rQ8jot42rdYhisrJj/C
EEOElY1gat7jOFTiRY9o1XwfipaKlIZE1R8LaIWMI06APGpefbpVAiZPW8B6+AN3VMq9DzBFOsFi
H8FwkD6UrMU7E1xT35IZUwWIpCr5CX2pbdfhF6T+v0NhNt+co3HRGgd7N9dUUF/plxRzUBymM7/u
vj5Na3RhaIbPrHIfRrpLbmlSfbBiwTlV1yIwZC+aefyyF7txn55846i6htNBkR7TnRPUYsWduzbP
YanFXzLUHayNLYdVO4v+8Q9U5NBNC3OfJJqEGU7RZA1VX3qRnnkbMrzjGkQuY90Z2oJhretHds7N
tuKGOHPyusE/ZafV1XkEz14HBw88N4Y/D5psE7t5akvDwG9U4kxvGKbBWMoDtwtlIZGqB6fELoTh
2Eb+LJpHKUqR7nX7FkXzDudq5iMq1aOeSBQy+POv9ycyZBDze0SBoYXcvCKX1gE0NFI4mX1FIrnG
sab8Qoy5Um2d5SxqQwRdForFi0B/MK7PMMn1PD5Wh1xCvDMPYHDQLGYB0Z9IXqazBlVoaUY0Ivxw
hqFOv7KsZWNIXAeBWwaH2ARP25Tl+rMSMOdnjQ07+Vi3Gf1nZ4f+EW+pr7Mh6c+kAAGcn94NgYqk
5saxSsc67NZ7TX94FMo2GyjWbF3GRuSIynfdD7c9Y5PUEWmNGuFc92FWjsX7Txw9sr1Lj9YGxO5x
DW+/cM+GFwNB2UflIBRKrMi09zMLYHYWoun7FVotkLXaBstID/SBMWQQG8h8zMcCbX2UOziBvkeA
E4F2Ype/2XNsB57rSU/v55d/t3E4iqLR2HZMZAsgplnHcSKZwWQZvvM3yYUjizebuAuV3Pmyv/2o
i2Dym+nF6ZPciVOTSav41y0pLXP0OQ5Wa8rCd3ZAsuAH2u/p4zXzNYLuGSMK5hHC7i0jfsKDblih
6gIwhtZ6mi3VSoB5xjLLpn2C1hSMiLRDmoi7xirBxbhFwy10Kda4IGPEQGK3qRRumDpKiy+HXxj4
BhjWk3/uDSpSeAB1MrDKNcy5bHCt9yyb2KKDdPpP2VWmxLtM/jxFMz+fBdqTN7iTGAJrkMi36+xT
TEJgCgern7wWT8S46QjuLDeZUxqCmFy3ccvSEMSNWlkbUw/g2yD/DtasQqVJf/B7qs2XgLP8lA/M
aCWzgJKdhrpApjAqX7GU4TUePFqYcF/Fw0zgoC2WM+kUvYN9vS2JLDJFzHNURZiwkjJFZP65f1X9
JvxVeWkADO1UAX6u17l/YFtEx1BW54+IEvCnHYSKfLOO4ljdoA5y/zQWbS0w+fSpS0tT2QwPRUEp
LduIQyt4ftkOXPmheSAC7jdOeuB4nU2QT8z+KzowDdL3vkQxJuuBvpsagXN8i0OrPNjLUk1hJAt4
9twsHlwdsmN0dcFJ8CqHJr4ynH4M44rn1fNt9i0iVCfqP9ZJbID7qoldgfySrC1PXtwYUQhJEAk9
1GxOb0iGygciaedhaNEjTDcFF82xShOMBa3WeCHGN/gjZnAT5buZ657dFje+O/MclncbPwLzZsmt
6M5JXGCDQEGZFk1V10EjYw4LbY1rTIpsxbm7TMsJMuW9xXXTxr3I3pDiySDCtv6WSGb5tSUf5i2S
61WxQ1NXJxBo6HbLjtfkFpglLt7whLUFldq3nELj+KGJ5tcBN5zHznKjBvyM3ori8Iauuu8JNilq
Rj4LVVyboZ8BMm50PAnNLNosprlfF8l9d5Mi3pgyEb37r3v3eOtrNJF01nPQjk3CFvh6Qh8fJ7H9
gKlt+z2HlKxnN3SWz7bigPN9JS2EIhrlhNKkOVMVA6Fzm+mqGwrcs1lPD7UVz4EwgeQkF/2nmBWy
jAl9bWogxnW3NsHyyESrVpOAOGe7j2+2vMfvpsH9d+vOG6P8nRFhVgP7Enl4B5p9UOrbEMJ8L5Oe
O8W5C63k/Cyal/laoaUx4pFbSx2ttStNVcBz8v2Lie3arWo5vqFaYISSb0qLAVwfmmIgvDG7HqbA
qZAeSoMHatEBuQzJOo2jxYMhWphsVL6Fn54ZCj5xVxhSWfOslBEY8PYmDKMtwxECF4u3WNQz/tsD
jaMuN0b5hw263zk1yB1hVSInXNR4TQFSg7TjjsKEwUu0uo7RsZpzcTe7BSaf90VSMzZyeavSlW8y
k7XH+0YTXSLNZr2QbSEFubM/qzXMGvYSsQ73QebKAQKnE41GLxDYMV9A5Q5fyIOXG2sSBQyC1RAN
+6bgeWtn2PlW0Hg7qt6lYpsFhbLgJATHIYQQdUnfWlCODML7bEGKeaqb5LZVLbyYIxerM8oWKGlQ
xuqCc2mA2UvPoyk6QF97WLcjt6p6yRMlRYg7Oofax4dHOQj7h7TeJ99hlmq83qnF9Q/hLvMM5tLQ
DhRlCVYcdc48uWyIT+PmavAETvRoP+0wC0I0+QN5t4Hjx6tceSs8mb3zfGgLBcwCLAk3VgAbHVRP
E4LyEphkbwZ+bj92JcH6+4h/iJ9CZIGmURey8R2IC+XCkxIjuL5uD//odXUWbgK/Zc4eBpDzUXqG
zTHT3Cfgb8tDoDvswRymymuEosLp7SX/XNHCQmbDH6qqrDCX9Z33Lk6TVOlanpyWsBoMMjQn6CZ2
4jj9H8lZr5athZzPXc7o2N+y9B54hwHNNFc3dquJ39/KcayARt1CKaudl4rz9r0gG9aR2oeBF1f2
YnKkZctvmSxs5Ke9HA8spwJK4+DJ3AGAqkLcuSrzscauIX6C1l3t8+QeA9x11La5xo+6ut3Ftnh3
cUHPmIaRmsBymJTRAtwxP/qE+mcx6rkeVzY9ws9hMxq7vrp6wiEmeTQm15yTn3BHvsKz2OBeVpG9
Yre/TggIDeXHOAGw9xZ8dEdnvtTRPQnstVYt6gaqTeQksA6iuE3mvRMhVNVskhKiFnevjpfoDnl5
gst6BO3p3fpbkgXP02hcJS2XDuUw4bPu6qGv0FBkoMS3r/klt8GupXk3ZoAcNcJEqQJsQpdCni4f
WeyfQ03d69WreopvqWxjCr0KxylwYlH4J/UDA0Pgol8vtfRjyrePJiZFG574CojEqPGeY3bNgkFG
rkfnnDRPb4pVUkll0rvl5K96QpynP8qigPZ0VIiO3VtUB0q1Mf4+gNcauG5p1h1IhYglDTs9Yov/
7+zT5cvrzknXHoDQFpjmfwMVbcfsybfitOW/agx6XLqY0OrGClu2FmL/CyEP5pP4sX8YaVyfFyGd
DHvsLbmXmGCCs+6w3j5SRexsr0AG1HmcPrAXrPuTCrLvex3KMob15pyGf5zamGtt8RXIktEe3+zx
R2GtxnVa+BXgOxK7xz2VmOyHhGWRvFa4nqkCJVqz4mkCOrSrzbMi67oL7iJyZyTQgZ7NImvGVH3/
DLAOejIRDmH7SWbQn4ykXi1Sg2ngviPX+ksXCL+RyAcFZ7cik2dXwotEWDmIZf3G5UqaYXyoaMZG
mndHgQJuIFrn2g9f/YjqUfYvxl2nlAEUjRGOXOoJKakp6IgGbQzWim69rGn4oel2gAqAEGSOyMtR
dWokdS/jq+XXlzQJ+PDYZ62KF4kNFHtwmsjYpHJ4w4UhwXGGuOUe0dokvGATQ/CVI2j8ZMlRo/k5
k2sXjGvBImv25Sxo7ohcSbfEJ0hBX3rbpywe7uXcu7JMNiU/DRpcC1ChF0bf8JQDZp4WvbWcAOhG
dIzGtNDBUFyyXgqjlp7e3Lz7fcQSoWByCea3O0/0BuGQbi/0YoW5GDtOH1Imv6bvyYm+USHnSnm3
23RsKPqDWnq1eh4y7Dr36CBSNCuBDBEvWnhtjWwqR3rADjT8jNtve0i8RO6imQAQteflH//ksXEO
pl20T8YBJH4SbPKawtZ8lVGM7DesfHMLRXJTp/4Dom+6wq0iRRlfpE8PG8CC0seCwuecGgJvghcG
L2kgbKCatQm4Q65OK+hNi+jpwKk3IjQnlQRehMyfkir77WNgSG4OuadHPykUu5ZBdWFlA2TNAVg6
2SF0MewJzl1c+WeUAUw6Nyv2sQF8IWvy7Yaaffnox2I2I0DUhGCtLfEtP9sR+8LpLDbJVkxUSYWp
kZs2Yuf0MlWqFjuqOLrG4ppk+i4qjIR54HeecGUErGiTDbPNJsW+mPLe0l2WoDQnk11Xlgile+NA
yUBQc7HCKKiGc+EjShwJhYX2fteicpYQMn3qTVicfeLB/0Ldu/59RbY/JWz4FJ1JBDpxKFF4Kj+7
PVZ3IzA70ZJRA9CUxjLIubYqHVTSuZ2C0LlC4ztHtYsKyx9vrHRTEN8gFRVght+5f3HjpWNH9iSq
9TBM6HvCTS34OgGg2AHmys+SBpW62IQXBSsXvT1QpljjugcUVuf2oA21CVuTokLYu0YCqcHJaZMq
/sodJrr8/DGACFsZL3G3/fmAKU27CW/kRNNhlYBOcIOinK8JWgjmWgqOyNXoACI72OMNGxTd/KlU
RaRIJ3mUOMsv1nlqFEm7pbar2Nx5fjWpnJ71g/qia9PP/sAHPeIbVSwKma+g6Cw7tqBdv7lUYBRW
jD+VgBXRdLqrzpHzktCzZgMc6C5pyO0yaOchfbjNOkvEAQoMTNI9Is0iFoUZ54JEL5Gm7LswlzB/
rvcawtCM2q+XMirtouLXcYiwSjy7WUPjnp9Ikm0LRVn14PwZoEtR3OxfHC4BwfurjSVPeO22WKHc
431zZjaDVnJSfE0AciDjIFcwU2E62oRkSV9GtZ1n9KQ1SMd35XVmTRfaaE4wuHaP1Co9SxXGMZd3
h/yxOCjeycKaXcUfqUzbNhccPAXXp6jd9+OVv93/FDb5W71x2uB4XPKR7FoRV+0l1e6AK77T6lBK
DDtwMb8HdLAJE03mBKushTGxI7MBAT011bNJlhlq7tTEwkIzh7mVqRkRplO4q6aE+v8Y+Bo2xA95
eEoEFwjmOmjOyBDR4ehvBaysYjjNDvfKIFrlCKYCRUjZtT518f8sp7YXhyTMVOFLMHz6aOWTh/Ox
VeQYdGcJLAsjxfmA48NYq1ves7C2fqclTXFBzDGLNYngJ32zts2+7+31937+DtschmUw4E0VCax6
+rgNR444WrgiYv8Dy7JunJ2o3b15yNEz5EBYDUWlwdgjdH8V5XMT0E2T0bGMXNewxXlxHrNwueLH
+EUIdXlXPClJrNpv5eUNXWXF4tifZ2qFjgJ4mN1jMc0dAqi0961k/NdkQMNZbwNH9X30r4CHz1V1
iOPvraQ/4657/nXg9NaJpLR9HW/IK0gw0O1bTlJcVDLPSw5PAgl7YP8iPeZQbtCywE2G0Y3YFHhJ
f8mZuGPrrTOGVhfWDyL0CMBO1rUZf/7rDD2PfBtPBs5lRfP0sxiwUDFphvDVqkSsVpeVHnit6yeY
FTm9KJwX1kFBS69LM4u++pcpGMF3cCqKlEVbZJxa9CohtOE7oAHxAAwXj+JuY3/T7pUDUnTkqQe7
zEX+eYmQRpcQnOE28Wx3G4TJ5uN/zRpmp0mCo6Nj9pLZPiVR2Tl58F+r7ItBnaWiwMQyTL6RA7xI
y3yw2zjFXn3N/7k+cXKTXdPAkaToAiARmqwj77krTjBGocOstsjeyo8wZ4Td8sbAeTGCu+fwTFge
PPoAZ+F19zoJS+BKjcMhKQC/yKEPwo68cdH3973mYYvWL+P7GfVE9bFe7yGmtUxmFTOdkRIa0DPC
Bk5mRP+Vno/k3462LJRHQeeszkYybwDItNjGvtg7sLS0sM7gxT2zhd7dTUxKvKqwx6RlBIgxJcjW
iDJMmH+DOMyGrgpLitk9Xvp5vEikPnbzUH9OZieYM6AnZiP68BTLpsm60BBQmcBQmvfV2NXB5gvq
QXMh3mY0jrJxCZGF++M80ngPqrTWEJLi6qzCfFyqcnJNvePmq7HxcF0rresubM1YqNPiDiARqHH0
mMl+u6uoc8Be47eWH1WTjiyMoQSaj2IFZit8KxYsRMuJJqPARwJuQWZMrse8LIlu9ErM0XDb39SL
aOCXs9qGUAwmjHxsFRtuPLcCqXKT//rSjpM8Fvk5u8FJmq0oHThEFCGusXBegtTY0Go7H6gE0tlR
ClOTqklh6c3TQF3O/bZxfs90tqJwWbK1ByLHqCd0XO0R9DmU6kR0y8+p6dK2/mQS6Po1+XX/fu4a
Fc4hmWSg7+ld2UTDoQoPDP7c2qsIoVzB8z17fdL/u8SfA9mpuUXbK+HoCLpbZu4UHErX/SvWs57S
Jbs1E9BMIhQKSXUQnJCGXkTgjCdmhp4BsTuw8AH42WCcbS/mPSUetxzs4XiwWkmiZXnmZhKy78/O
3+/eE92nTfYYqxDCdyOMDjuuvK1v2YURnL+WY+So9rHcTToMiI1X4bOo00lgKYxpjcpLCsU9KFoo
zqPK+A9hpp/tdY5EemTmXGbvozWELfRVzsBR1niNwg0J2Db7+zii3EPvc+kXxjJa4K6Cfnwhx1y3
TbzDlVJMv9dPn360iaDLOOpj3sIsy2pOrzvlOj9D6rSfkl/YwlB01+4zOgWvkI7WXAlACdlosmTy
Sm9v1QiXnCfP+7eXd3VLo32qn7MVunVAtxDC0mGavTCrcoKpF8BGEAIiqSbEMsoQbD/0xMebxVfv
2RRZNwcg3bUnArn8kZ9NIXQSJ5ZHn6b/mI/JHEkIPKtTNq2DfUfFfDV8JYJqvz/KnGyyLys+atmq
Wz573HrXFwcsUjkV9GafzkNOozwET8N+aPBK1HuAhEX5gJ1Vc2hcjqr7ozEckJa0hmyCfFfskLzZ
X6qvt/g/I50e4wzxJwHLvOSZTd3gX8INeA4lluo5e09fA6ICiBpnOPBfLfl2TpQTbUQX2EQRXrEO
iX8vNCr1zcg+jqoKqNbf4fsajkeaVwcAHjPQCXsFDVe++ymFOq7/IHJ9NG6oCMOlJMSF0CDG1cMb
gJqL6Dyxxtt5HVFykcx8JLeqVTTU+wxE1zsTkdzf/fXAL3EopZIrhNbEL3/S5f0+O2P/836+00gH
rz5jQ10hXB3kfUTltbsMkAakhx+J4DitrKt5tPaWVW4QmEQaXNWq425qxUzc7ODOOWQPXcV6SwYn
uodSWHfkePa7wt+bHYO6IRQOttRKoaCuB/J7O8gkAzMvI8vloX6FK1WHlbdCexGzgOsrDkZZaT8e
8jUr9bWrRByu387TXOJsx2RVeUZI765uL+H9as09Z9Wnw3wEluzcJuuwNwt97tY0a0g1tiTV7eZ6
FIDTEa3qnwG6Y9eIKkc3krR7sNKd/wyshLOv/PTVfd5kXZ+og+l5W43BjaorunPeK043wEBsokOx
3nrd23b0W46tvjtThSjCXDRYBxrEakCoKgJKOxApW2jmDxkRGl2BmxqCuhKloZpyV5uUDASTMnQt
QHcYpjo3BTZ5BpUMS4ifSU/RcEQ+jlp+whVDyhUirD+76cd3pRq1LKi4Y7qP7X8itNTMZhB9R8tW
o137eOantO6u8VBSlwRyFGueorG7pjjxjlqz7Njubrx1I6Tea3UBZGY5qtHZ31Uw1fLmZujZ9hZj
x5U9FbBUE/0QB5EueHZR1g2bMU3IzUZ/qXq8OrgioCBWvLpHiKtZYfEutUHskbpxW/6ZBpk0i1uC
nF2UUDIEm8o03yWFSqs+vvHAJGrUuuBHui8RdA97/cf9uU1uobFIiKqjQiBH3kAgVUnB1KlaGAq3
xn/BKsu/UcK+Xlj162BSBZYDDmU9v9xfAtyeoQw1UsXyoQUm47e8LE1fW5xhZ4TXDaaITPlinYfA
lG2m0VGcDE3rhFYQeeG+SDqivZAGyz6HI/p2dUsHXf5D9QxaeLqu4a35MAlDuj+C4Ly9RldGYerB
PcFDNUN/Qgp/exZ2b0aGWvIQ8t24q0dnqT0PHEhQTbX0VMkTDo7oIM1X1RpcS2GcM7Nt02kR0yBi
TS4456fuybaDwac+zxTB7D1wqsEhAMJo3fAR5hAckkz5f5uFU2oc3iboit+WrEt7DJ+ct7m0LihV
LRAZGteaQV4lzDVvTUY0o2meFF0qMCT6VPsiZSXFbTsloSBHXuBqN1fqVYa7J0+PywSyxPqlCRRG
MyfFTPn/UbvOv4uQEfH9nCOQWWjByVxwfWcB5iy7biQOfhDnMZdDUeGl+AzXPg3Y/9Q45fky67wH
fc3NwUGYTNPt9/UJMavkrBWjvvI50vY+QrcmVtsnWMEjtksce0CoVUgDMG39cI1N5F9HX+EPQWYU
TzRzFIPrZvSXrq2OUlNvt6U3Z0B6WqqznIXw4AK9uxPCHMVkx6CVElMV/kjibqRgrYaf5PzhSFjL
As+zLmLLWWsWfQxRslBzByT16wkjBcnJPxLqm+fevesFhz1ZujnFQCo3D6QE34PS/+PhdRUvNQrT
ggNCCPl0wo2mLswJYjclCGX3cA94qUJAWBXyGQ5+J445qheew0bqThLHd2o+SeuHj4QwyxRtK9Gw
MaVwlzi4R7ovE7JKoTvQx2ps1G1yUujU+Apa+FJvdUT11B5ZdTindi4dDBLnmb0sgBo8DkFJC44s
P0c0POwnKKJ0+wDcKfEuMMvfynLaPPWW4eIHxCzR2tFcG5gcDGiBnEWoYb/n5jBBzJ+iSCrfulaY
AYddbL4hTyArA/F/WtVxkMIzqrsuQC2TgD45KC+k1Q08UeZtkvSwLxfCnm0BFQinoPGaTM7mNTo2
fgAAvRd5PRSdJE92iVRu4NfkvRrF11+8zz5x7Rl/f+Jdcg3xijMbj2/BILG23jA+wk5rg2PfxYyE
DWFK3esXu79EhoPnpuEYqpNbasiNODOaqLZsKs6+et9MHMH0ljG5z2AtYQxNwRAdPPLfvIHgoyh0
3u/Wh/Eipmt43NLC9gqtZHaOsYDS8daQ+xH3DvTh6SaEQNdRfvAsgL9Mlyzqgt9fo8EXgqrTCgFm
kVbxjVR36NCtY7Nm5U5SHl2xW0VdItQSNZvocBlehA6PoxQZWW9sBgGQJVZRxzyrztU0Eq78qaSS
pkRV8vp0TbRx99aaeQzEao83NTkScVPHoQWzHYPEcNWYbjWa2XX/M91y7QqbSGEAEI3paPnepiFs
gQNqCeX474WJsM6aGdawq9LLLKlbGdMCgYnUKnIP1nhdysZp5GptVxh0UNUltUwbLsRK7XjXkrA6
sk0M61Vv3Bmv8LAT6lRIGhRpFJbuQNSaXPabX9kXcNEWx0fFRILiK6P6hF489muRi4H1IWgjmGqN
fTVyyUrIfQtkhOPfbrfYxMRrBTBW1GTi3H8k1Fh1OrfeL39GXvl/cf3EJ1Jcx6LM1BM+xOm/XGBN
d3fVWaoXJf0cOY7Sr1gKcZnXp6zJmX0E1ci9CzYTi2K9A3xef8I1ScN634ozzKarS4D67ZnX1xfc
D2dZqY978tjQ2YlaXdGmHJZ0DRrsXnJbuR5Zf6y0M86Xc1Qt+NX19zwjBLHaau/C9IFTG3fl0rlw
haAJDUuXgDGQuGRkfTkiLH6djEIK5Tmc0WNCKDe/DLwVLF5s2YDyPQw+Rla2vT1s0NoXNK+FTJHy
SBvzssednHy909pbm33pyJYRWTqvnjnFCorh0e7PDAN8bRoFwpnR1DcxGnb6jfQA3+tDQ1Y/woo9
Bf3nZDpAJ0YAK7u4wtiem/Ax0/hRMtq471MJznkJR9zK2aCb4FfRylMnP80RSM/6EWsyNtbMSo/L
jgeE5CjybDE7lQSp7u/mW2AvBug0Y2SWbyi9w4dKhj5uHt1ENjBKMQIMYBlTEPS3rRvCp68691qt
EXY8OfaTcmF8jkJvnZ2qjWMa82ccvynPhqYX5tW8IEGTZM1uEmjGc4RLZeTASP3R6vdWdUzw+WUP
trkjq00BQXbG8ojDFVLE9I5ohJuKQb9OXhjo6ZpdN+3j5WnqiKQh4jpEfvabhfPMBYHDoan06wwc
Mr0qafuL4c+ubeHQzzPRPP/mvSzY1mz6fgDuJ0H5si1P5SHbPO/bH9ojOHNjkDnvRTKr9O0uJXMP
UgnDCqz0cMkPZluQnQZGWJvgYc7LppTUzYQ/IFBTHGgoOYUj3GFyxy2EsHK14AidzuXjVugv1UOr
H8mxTGGW+MLipdHmeb2IUBiI+B52JWQj72Jj+fRvCly2VImDaA9ol1RJYA0fKThq06xecU+ECuAn
foAq546bg6t2LFFhasI4JHfd1ENsd21Pzs/uzC5ZSfucOgfc1evAOnHuRyhgqzCJtQobMGJ8sgKY
9ceBYn0icZL46KLzI4AipO6QxII/APXHyK6P4BwXjvuJ3luqyZIndDsKP2OustzQqbLhfgpReSVY
iavZl6SHgZ5n2BnLQn0NLWTCrIT6sDxGajkbx73boDNntmK2HwOZ+CVnutRDBarTeGJJPhA6l+FO
g2URtXymBQueKhqsUwHi62/bQaVWet3Ksw+hlxkdivY72K+Vc/wu1ihYAfMeBRv5zi7NgQHagj70
Z6i55l416hFSxKX9CUpgyN7Xs025kiHGU02KPEuIs/j9m0ky8J7oadxJJYa8XojA+E1U6qk2Qyss
dRpUTRsrjH/wRcZvm0u7iBCeoPBLYularKu+rUJ54LIB0hNMwgQ0HG+3cvQ9uW3O7Z7Rj7SUhDWO
unNsHaqTgDZ5Hf4YUUlxZMGP3ni8qhi0uUue1nvbNTKQhNkV01MiJGVF9hnOopiv6GsP9rmQDuku
0D7v2sGKq8ur7p3piXWPtiSAlwFZvkSsEHbG96BUlku4L7GGtIP9oIJDtqqz5LG+0jVR+ycazt97
3xPeUIEJactFqnJiy+Nhfhx/Pn2qnd423vz2YU18S7HueTSr6hfoCrFaHGXYrLnSZ9f5LNNsfdRf
wjJGkU92pCF+niwuuwUPp3dYwI+Sht1owjA5vFkvrHa8Q2722PjezIfshBkpf5QJA4muAZveDDTu
7RD+MApRfckuZZIXtIS52bGZc7ViJt2pHjZ/pDemtg35pdOgvVDGFAHXSg0zMMw9y0wLYlVqwYhO
3CU3H/meOHbDuDgZaUEt1pr0axxdaY+zY3PettDvqvMaYLlqd+9nkulKEJxUAG515mrF4QMQ/PH6
M/5/JZ713Kj0niSgAzWa9hS6qoeV5iQ1g69aeR2ASFOBmL9V/eZz9VoMpZDJSsDX2XrsqzhHWc4r
sTAs+23NCeO2sAWUhTp8GrtmbVphvcEUvNKhAqaIhOERxaTWXbkn7p+ZV7WTxgNVQ0cw+71COUx3
1HKzWkaLpqDEEBbxvOS0SZPiWivJV0jM6FSfIXz9FtEUItFsPNf66XOK5IrW6Q4ILCsktvmqLo3o
C+29qbtkHNl0GuXfI0j/ZL0xvhQoGbcaYop9FoovsNGksgBUuhyC1H0cdCxciO8sFfFX7enOefqr
MBsiX8xg+YhRFbeNUJXTuK/W2MPbGdjaC08UyYuGvsjq5uD+Pks7pXWsWVO2iyoCkCh9JdcIbe6e
CoFRJl6/15J2GHD4Mu3grWCZTlEiebZbMtpbfkcLwgiu3yzih0xw0LjzZvSHCsBdEMRJxF+Q3buV
Med1UjE1Hd7ArHsJRteg9+R2mR5cb//ZKoP/NMDm5ABFIibEDqH4aSy3Cdkxk5wtOiMhlnTLdBpl
F0VSR8ZJjMbu2GbfcvBbgRKTTLECW2iJGgnKWWyr/av7vdmWwRyTBJoQmJNduTe+YhiJTTiyzRDh
gRNgU/sxJcNf3US6hKt7bIjZ7HlrnOXHnpy846rgGSKQnBRhXXUQxo538UFucnvhcY/YhL/rqtco
zBz/olEj8KFTacScHBi6Z7jcOh541ME9dL/6kZXfetDlushUXRjrTl8xBCwihZQrq2ubFRRNYTub
214n+PjO1QjWRTuV+OVCNYHW2ejwn/N0nZHX+bJ0NuKH+umg/RoTKFFtOQPBiWZL1cbQM55FXB5c
SiSmKAMf9DutjX/Ek3c95H1PGBJ683J1skNqLFZwtzC6kQw9AVuLZSYlGf+cHOVgutaxLFFogFmW
8HoBqLU9qZqcmdvYARswWiBX1KYfDaWwREzXAYxjhhVDinGvgYX7TyMU0vZtcJiN7cLn8YPXofzX
EomVld4OOh0obf52ug+j9fgO2wUmekMAwrCYkm60iMM0V5p+1fFE86QAxRCuRCvx0d60V83DFJjj
KcuUtdtArXh3g85N10YgKa7pBkEnhd0CJNTOWcboiLP3tG3sahTm79iMIj2tX3JQ2cAnBA/4CKoU
NRXDqQQ5Kp9g0rTyDWxHThFfJBI2GSO6wQHQ5YVahEyVUxw6pGlt4Vz6uU/owmNSlfgIsoLd9A71
nzxBIp25Jg5Kcm6TkwdlMLG8TuaoA3zmI/YjXwUhDJzDfNYApkED2jDXCrDu2zQXNY+tXCVqot12
HkdOWcgo+dsv8xwAf6VdbezXW19XMCgs6dg6aBNeba6oASqpcRREwS4Y8p3+a/vRh7qA4MF+1/K+
+fajrc0HaYP+Ie1nmD0ds+Pr4wRyeNJ0fP2gq/Ivuj/7C0oLizmh7f8wKsqIIzXwyK1m4EU57Ikd
3hYzvZqxyp/2JoPC+2C+itT0CuZrvF989/p98OhPbn72+oqLy3rrj82uOVq/6AbKTL9ug5E7xtLZ
Dlk8FC93OiPpKtNfzNRrBClRaFrFqyrV2Z6kotwXqJ0vHbV39klOV0kFhlxQ74xIsz0xxeyfFvwe
W7pw+RZ7877QhXMD61Z7/wiS9/Xc/g9ZF/pxSQ7WcaVIK3kvk6f+2MauTK8HlTZXoGfMsUPSqAlJ
LoWNusx560kOdEbVS5x1bX78kab7zcyd9ON1OCtVPj5QOo6YmOhGPkr1z+yTljhyYhzF4l3I8Th6
Q5yNLXJxIUXVaxZTG+5FFrTDEGJT1Zls7riIH6qAr2NU/srXHQqOnyH+t5Sy2WJWwrhSdUMvWuYC
ou/bJiIgNzfK3+JUg3EDvV2mzMXK7qiAWwcxxcC425pOdWne0+Hc7Rdb/wCdZZM8BVnY67tZ1oT5
KXvH1EUZj7UECPR/EfDHKenJFJlIoa5bWYM9jWYZRpRmSkI8qHS9H0ga+kGKBdLZZXINKGZzG9iG
8UGaQxBiK/WZHu1OHzNZShspw2pxSVpgRgXailON7nJTWLHqgBs4L69Y80SUE2CWJZtSOf/iwu9v
yBe7hyEc4p7GgufYnDvFbog59MTSOH9OpY62v9y2Iq678sB5pl/IHNOkrz8cVkolVcC8Hn/L3zgW
PN92i9rEiwNB/GqwVEFt61eKnitjQllGVMb589V04GRqqtj8wuFyIzF4A8StYBhLMj8pwfqTLsm9
HvjBGhkzath2AjED1g0FZkWxRPJE7gfTzOb+XVNYTtU/jzC1K6TsOoX4+BiefgIpCNoc3V9cdUF3
E5OPAEPi3wZcXFWivyF8XGsejsUYDG3tsk7zEtitkB7e4vqwAUl7vGnHRURknZzu8CeNlZGoJnDe
rit+qvy1sVQUkSLbLfoAp1jnoD7XShf/8SOcuzHCAo5XBgt20ehV7osHjwuayHmDrIO3aCLxZ7iA
01ukC1mQOnahtV4iixIYPozfu1I1We3H6psZt0WQgU7YPMOb+Qrtk8xjsQChJrr5OK9zyOBLVFqJ
+UsUf9wbOiZMnCDBSiz5FVU5RVEVl7ApKgvEwOv19Tb1RUdMcUYdakrLByrsSGoyCP4/ShqNKOMM
8gx4qm050vQfj+t7YJvBAyvvNwPDPVgmH8/TYVMbKG42vUI6DvSOFftrEG1gi3gBVGNnxrtWfpYI
6tMb1haMFcbr1MF7jaQV6XLObx4eguCrskSq7ja4KeBmjSoSfZv3a2ule3A+g1RXM7DA1D79M7Mu
BZzBXdZK0m/9c1AJkxWxFshhgQBiDG1ePEFZAuB8uyFOx2G5cL4z3pH+bQyI2NiUHbIFq0pIZ5O4
kCHJhxS3dfwsgEp8dCsfdqDt2k+yVsoXd8hHwzOtlVi4jn2rzks9BhDllLX0wgmc0121aIcc603Y
R70w27CBmninKsshF2W87UGe1EwYHkKsFUURks/ooNd+tTB2loQQoMEDGPgRhRkBtTvopGiseeGX
sU3n9u4SxP5XtBn8x4hDsq08bc4YZV7YU6JloyeQbcFxLbee7H5XSMgqzTpNMBh22C0c9zrNIZwp
5xUOlJT66gNHD2k4Sn/o8MOWL0SM1ETWdbQ1qPhERFHqc8r5E9HSiR0dKqTm5VZPrXwkL90ADTVt
ZHCXDWtR4yfIesd/SxKzhY7uBgmeXSw9wjH8CP3tCloQRcK7AAl9zIWia+64Pi6QaYRO/oP3o8a4
UMTlkoqNdwrlpxX89AY7K4jYkLYWUz5zj/3X14Ms1yABRpWcmnQCY1xtoe270BiAcAHMmbT6mEJV
enuLh5K5k+b3V/oKH57e0z5nBA8aCF5nX11HI25kXFF1tH7ZzmRdzC6qXkU/nLsBaPv/NII+j+lB
O3H7trwcdckpcJoXvTKHyXM3/XI/8iq6wBxRTna/ZwqqBL9QeV/ts/GNcRbJWwEgx8BZNbo61nbk
FFPlE4QKZZBCDS+tQHTkKwt/yBaGmZWB7tBFpYfAFbr+cLfFA6qGMfBSH+2TYc1HfKTdztv6V9yV
AzzTXoXVhm6Ar3NRso0JyGUXmurOJ7YagNexMSgJu9gF36QaDy9kPYC0iNuchVZ2r+8JF/8Z6PTa
caUaZgnCUn269mpyZcKCi7gNg7bK59FcOFrj37hWSP2LdmYtkUQgeYEcqFGscB/kNFSncU64SwXg
QeY3VUY74uL35+Qihg110i+SWSkRxp+zPrUOv9gXkyT+v6RdrcstSs2yRMkfZ9xFfonXhYoD7ONH
brUsT6EKvtFfsxe3Ktv0XqTc0XmN1iPT1SmQhz23VuaVumAYQrNibakLjXLKH+cgwPA3pXQNJggf
fYV/5LLJPv1LDMQ0cjiFpKDv20Ta0lZhapB9+EEKeMQ0Aqlx1hUZ08zR3wxuVnfVOaN4x4NyhFCi
xsHO5vwZk4z4UZrS1Xz6QrnayuZuY/3Gxk3nepFNlWTa9UMPM+2I3GxCPEdWrAG+hALaxoNTmR4b
IOtoSMtuvAANx88yrfqJwqxXVeH65xPT7z7mj4d3sDXzQ2RHd3br/bj/bx+McdFCFhjFKUvTTgkM
+7QzSw7+SIFAlnt89UwVX9wZ5WiNu6ZZzvMghaI5rUi8hgEjPm66t/8YWfOZZM8J2u3fFS9Jew9V
hKIcRI2A0MDTkLifqzESMYymHpLBq0grUk2f1r8YPvqqW0JV0Kgff9nB22rNtT3d9yvUmcmog6xO
tENWvEh7jfBu/bYjcU2uzfGDOFJqLv4HGMo8djW7vZuBkUa5H9n8sLDefxwNiAm/VJPrdK293kC2
RmFEHe1ZXVHa2z/UH/ch6c3H4nmRsT3sWmL9cmTBil4VqtUJ+HtUeS0oQddRyctRtZqH0ScCJGdM
0oLGXdZML1yB91BKfeCxFRsTiMvlKXQ7Zx+xETtFtfg8RyHHh3iDoRZyrYGHnoUy3wQ0f3eqWXXw
Z4tXuv7LIpH07pSw3z1fCe/K37X754fkiSTb9+8cVmet/lw804CTc+HGAcobPbnTBNofeLseDCp1
D/NQlKwWRafhG7agLClpXzThfusDbmEbky6f+2IyXOab+sBvkFAOLr+8cP31gLtxOqWig2DO2H6D
c+xsOWQhpLHSGMoH1JaiH0LRFw69gB9F8tdFa86IYCJ2+cSI2f7R/d/ezS/B7U23dgKWlePrbqnQ
XJqnqh/AdZmGBUEDMczDFSGCf704gYWcg/uUaj1K+Rwz/r0ZNj8EV2zNd6TrWrhVlRSx0DsMy5sB
vIpijk9VSIpv+a/g6TTV7ZfK45wfk0Nj9J8JKgzPpKi69tyUFFTOnc2Gcy2AKWnRT6J9w3mBzasg
+z9vzj1E2Gl4Du0oShfBQBPCnc/Gi7+t3WPdRWXKljU7IKi6DNpqDxeg5syHQ+t5vtjNlt/+lHHJ
5xOHs93IlIDTePSUZgjorKY+WXSHRah/2tl7j4WYIpqTN4Z95pckmfTUnHmWE/mt2RsoBJQWaFZB
Uyb2/X45iQf/LNnqFW+lCgjHXw0eiaWbFVBv8lyUOCkEG6pR4mTXHDbGm4r9LyHC/RFcoR6n/L9P
d7wFu0/YILmWoWDeetxzeS7DdIbJi4JqsFzf0nis2nFZ6KtEBS+sYHR7CHsMza+z8Rsb2vqPaom2
pJpCu65q0kDttFA7jAsRb9U6dUVrUgg7pR6O05M/fW1d+2bgniIDQGQXSpudyymXFCnL2oagHhn0
ypj17rVcWNMHZzEJHvY5asucTsG1jWNxpJsCJ9Yq1flm6gLS3YKeejFaKZ2KSaeJ3HR3+daKSJZs
WxWiEN48AfjD2ISoyESxyAz8wxgBrUH3z3fiJxtPHuCujTc6F9yW6LxV8ng4Oh7O82YxKR09izrS
hrqeIAYptNI9YivjxYs8GBOHNG+L3pLIIHUxpbeGsx4ESwZYFKCV9C1MAch2r9ZI/9iSo3Qb6H6q
Blb5uRqYrYwkyQGfl7cFamxPWz0qYPhmQqkpoP2E6ttAQ7xLI4sKBfXjOR/pJcW/Rxdbk7mbS8oW
IWoPii+v71Tz44kUp3CJNHKfgQ9OAhHynLSgaNETeBdvKJjuwvvG6JCtQNzU1tt+HviIdmB8ioNs
BjD9VNn2NjUrbpLkQMCsJD2Fya+UK5lP6wyRz0m4EAzX49nk0B6IpsPnfNgGiMr3q2/uOtEiFll4
IRG36tSe/U4TD7po76MtGec8gGZ2MxRarqIttsJ9tR9RNWTIMGGoMh1oXV39LPgqkRYkzMrFC9hV
sSjLMomraWQFS4676ZgH+zPYLe9D9uQTp/VqBSP6ChXf+hUM+3GW1QWNh0UmqLG7EUBXbLnN9OV8
AjujSrinumCrhGqO7WTlaIX+yTmXVSn3Oo3ieo3WjifCC9/Z/NkVVNblWZspSlXoyEpoD0aaKwXW
pN8k1ZFz5oetCIZpoi3/PGnayjcyiAXYoZXKuN7eldC0LI9jlMe3whJSTgzdvDvPfID7GEaK23dr
jgFTeA+oDtyLj9vupFvsIRScXTxahD6Xhbs/GK4AzK8zrLohfNdDAIndivTwKKLDML3iabsl8Fmo
84gCodL+uhz1wYMw9AlUcunVelNGjpKCjhM8CtYX4GthbzBjSNGZ8FucrKwqjLXRLI4xsTvOrbvp
tdFvzwS9jZU4iyYVOSXJbOb5/0HWCZRFjFY63x4jOypNOASgILc/PU9kSf0klmTNG4/Me+hw363Y
uU8e/afCrBZ+uEbz1e6cv5rWi9MNrZ1gUP60rs99fZcJnK0V0rcBEJj0eBENYCKGb6P88H9xFRI2
bWoNDiwHtM1kCdSZ8fOO15cmkol3QFIHK5Nn/SRL8HST/1dXwYNwj9QzOIlpnd1ASwEWCBhx6+Pk
bkjau20xHYu0EVG+8dl5ZV76LjrCgVM8jA2bIBPjoi0BmvK0BKAzFer7zHDCPABVntosEl09KY67
UCzhzsFnoIr9ATJ4ZuEUi2D5I2xqjPWEx3zhwj5mgudEG70rBlBTGev2SNOuSWq1ktbd9IfVgzn9
WCeOOApTLmovBxGH1fvd/Wm8BtCNFCnOV2vfPYEOPOdX0ZQc0EUhehMhx9CNlC3wage9aWIgkJQ2
4YyxbbncXpYyzec2AoIftQKng1BCSoSguLlpt9vKXtMkZOiCuDHN7bBkeTgbAglnGrRZYnjHbmI3
czCR8JCNCsRPZgdskTcCgBvaOjcvhzbsLjOTxTr5nxgFfmmC7oKloxIVK6pAvXv4GtrZnfpKnrga
QyNCJ52PGlciWUC4IPN7LmC76sfzKZsqjvHDc3ItXMQWpuqJ+lKjKRcOliY8yUHdL4wXvRlWw6Nn
5rux4Pc23bpYu1Um8ICAx1F3CpP4InpSlDVJ+nIduROIvo1jFUIVWsM6yVXaUiFs1mIA5gl6GTeJ
fBt7fhXalMBYayB3ldt6rmFmbDVrlsNrEQaz2J1KwmEiZ7iBUsXaBKcuXRTL9rAt4t/xiim4pHfS
sYVGS10Har2woLJ/P/ZHOoUPiEUSramnHjxdtGbWNOIWp6WUsZedWs/0dEVbv3cZgmRU/jntaUgX
KUJRKRDosK7AIexVwD7rWRio6UpVgQ2wWmNG4Wr+PkfV+54UIhDOADXw5jvGKZlFOIApglP4yU63
iL4Lm6v1POkadEbCzo1UowAwuS0jjGu5n5n17nJYwHiEZKAydn67q2bkEu7bWRlCRtAl4VChvWGz
ohQoNFdi+xVovH9+aM592coEU9mfJaMr3UHJu36ISWpFIUXZlL1EyZ7ROK5XrWlreJjTBTLyPvTj
L4UXNtJ5NiM3xZW5e/j5JrEYEgLVetUNhnnDnYkHBPeDC0IbJwNjxIryIoZcFVzMYwn4yDfT2YbN
9F2ogZwx4e3/olozT+PhB05zDE/z7R6Wzm3pUXCpZFBoghdtLVrKwOG580gwVSrDHlW/FugEF/De
eTlfcYA5AOGaTUhzu+9X0XFg/4YB6aXnm93ywkos9pPZezQG92p2zUQ4mp15AqUbADd1/gMXyBFM
gtrqZnYzvHcHXtReiMSnudfzFXD7999gmJkdV3uFuCZtDp5zMhTxA78X4dfnjthec+jT+lY3uiUl
HBzt34lACDMIbu9CefIbQqum/C+m3I1LKEy+6pzyBkTgYyN741zBwr6QAek9WvKdtN2S9vUxDsFG
sz0asc52s+CBiWhYfDPizevGuvtoFiZbrslq84H18qFi7+sFlhY4Th/JGVuCx1SFiiY5XekUdsi9
5UqWJxZmod7ttTWmSErYKlWL4xz0CkoGqdIk+1unlmtkPLm3ospWJXTY28i0dKwLY9IQfgJn1Mwv
tHoiyWYc1/ytP/n7+bYv3xYaRlr4Vm4Tk008p+SucBd8U1+jsHPkgZUKC2V/2khzv2ATO8kFvfLT
haLLX4DHywp9xQTw9ePPtLApimIfV5DiiGnfzXfHkFz68Sg/J6TTZ4CC3u11fha+tS18g5OzbUy8
BOa0zAYH6MMTSWldbHFMbJlwb7PyHgmFtHPc/qOZXm6KIuKy2HJoNA7CSuaPlIYazfmbXdxScC8/
Seu9QK65yqrlTSX3m+fS/BUAvegYDUPxwrs3c6hXOijf+wXkDDMd5vJivU7Pjycz/9dkjTUcnYHB
tOjjHV22n0VC4cxiEnrpIyKobmfw5y6M1HclhSki1pGO5ua06URnEmPz4l/XhtS7aV/8qjjJfric
PzUluCRvmEG7RNY+9dlRpW3p+M1ucP/UOLtR9wtFhwEqD+CK1KbfCo/sVHvZrVbozGPM7+yC6X0Y
4SlvWUPOJ4rX/LsSwwGU+PbSDSd/DeRQvggbS8DSi/gD1ouXi1orRLsKaunTWFwQZA1T8WI5VyjD
LHtKQ1QeOyTzc/0qg9+oeqSgJTheMJ8tR227USWabiWtmvOLqlWJXdGT0owYXQcg7AyejvshmqZb
sQzcNjgQD8yTi1SFVtV53fHlX60BQ6lgxKeaVzrsDv48qTSDdaVdhpRlZRqbY64C0j0WmUwzK19F
gsWW1CLfoPbSibZ/9rTrpH49vDEwAnlgYPkt2wtS0QB1IB2TonI0FuEdbCPl9WLaFIvsCmoAhjFr
dPoMGfkSw2d8a0bMLKzxs2UJYCFQJgySdyX0NE8vD0PzLdmjdEG7dlFbet3hw4CRaWA3eee0bKg+
2gUJcLSPoYsp7Z//2+QgysHdxdpE9ouyeuTqyOkDjcMDxVoyLvnqGpjFvNezs+UdfCwLqn1o3vxh
UKXihOOh6X9fss3POFHK6f1UswEXFp+6EyrCMHcp/9ues2VL3Zng2w0bDDuVHe/uru3ipE0c+y6S
13qU/mt2LI72nyW6FeHYJj4xmdAFBBKtu/nq27OelCNm9zZ+uK+nUmJ5ZFOSHkshbvm59LT52TaU
wbbDZlncLEV6xYrgnZOe/+pqMuR9kRlcNjtYGc4vmYyqtDRckQCttXY5YZoKIbpFhymGBTHk728t
oJQk/6ZsDVC/MrXYT4/ALlcqJ4jbx1ZwwzTyhsPPBr8hhz7Xjp8/s8xW8qq3GBjgitOU06b+8FIE
guVrg43EZv1NX4Ko/fTO9doVdzSA0j0G7Sxk3ugBeBQgLsPJykWIKNiDdk1SDVxhP0wuGLAUdHe9
IWvLvsMggUHbspeBBCKkoP4KOJjKpL6qiN+TW787mp0bKuVgZLSfvL/eL7F1mrpFVAgSq6gTuEyr
aEhSy6GFnDnDCyorgj1bzUGFqdAqI9GXr2M2wSd7ttk6CTg3dq5Puw8vKBQ684W23j0nf+hTUo+u
5+9AjesTOJGhy3S5sdDBVfDvxZXE+mT65d3S8S5svIJi7cr8ry5saZbW8AJjNAXzU3BOBV8m1FV3
b1iGvYTti8LkvN+uWd0R5WOWLhAndi3snrddOMvx5+zOzjUpBekR5OkH2+N0eqfDGHSZYVFoi+Or
+vwxyKiiZgi2VaodC8qs6nLmQDrJVTOCStTou3RnG8GGgGS7M8I9mfkWFODbO09Lk2B0R4fC83B+
sHZ/inRcjw0Vs3x4ZmJfcV/sr07SgHKO3CnE66Wmh4TnLgdwF6QUMR80coPIU/OADDLbup67rI7V
YxAYSFAlrb588bc/1hNvWgHGykn2NSUWcyGx2XdO35qDTaCVgsJwpOfoI9Wx5SBOogl/NVAL8epG
16ISqaxdQCEm556k15CujEh7YB5MPIv0GTWAsmD6626GEbP+7DRizpVZMjjFCkhxy143Fy51+rzy
a8vL85d4a3VQ02YXPzWv2PCm2isAUedk7kvDmBhjYHvQR3zozxbe2P/j7E22fYZAzx1Oo/uXz/in
s88Ym088985ZC7ToQ6kiXEhZaYvXCiFh4/jUxSztNxtnwNTpiTo/oXgJnp6ptqoMkLZXi7MZPuxA
oGjF18BVcLkoetuXA0fnl5gWdOikhFZGUjHm0QLOPV8RvL2j4H1pFiBZdibNHGJtUtjqp+0/rMnq
IF7SoPWBzq5OqKXEWfs/NVey282exRtBzvJYCixk9pIRsi0pNLsACkTE1r/ShxxggUq4ZYwD02wF
u24yIrYc7RnewNxcGWnGnRLV1RHPbc0VLd7dyikIU1BXrnS9wCw5fkaU68x8fWRx4//ZB5wbMT8H
TOIICM9XqzTEB8ibZehGaAkx+AE2syE5bEOiTnFje+A9Gz+IS4QPrFDEI7ViOipSWuvxXbLDUH8b
F+NdePVQOaP+PzjbjdePrwNfEQaZo7x7j4qjfnzKH4uHW774Ag5rsx+m18WptedarJFH7oqYoAtE
gGIrsGmic0KepqIjYCTwDFJgWSXrbWTraTGr0mfuW6BP2nfcc1Ymnc5T9Xb/xU7p0jZTE4GaGDB2
TlVIquX3nDxqoSCI6/1TG4XAoQ0CrFnzJqkiTbHvTbLxc+cm2VndgS7L+rG3geoujvjMUaBN9zMJ
wIyXkTYnUK5jTrNum2EXzTdPha/VyLLHO62Hzrg1xQdWCYH8/GtwWHaj3UILST3AlpwqmoXNiJgn
Sl2YpKQjoVEtfoy3E3j9H86SH+WLqBcP1Z5tBtxUa7xp5E9FmYZFGJ29JZpNNUftgQuL405BAoEG
woJIs44cj/gSCNaXQ+/IEO3uX/0Q3VReXYb5KP2B4Fw1F8grTQPjbGXzx0UnhTuqlsQEvbiiSwzR
H3cdD408dd1/t4AZnFQ9/Cra72QtNoI71jazunxDdWcF58sIGHXBHFpjb/y00X93cGKCXn4uj7bZ
t6YTva4jxjwv+d41CRS/wuSA3mAklNViZzJtgBVednDAKngQ74+rvXA/Za2YwGw3Fjd27VNajCUO
2FM/rN4e7UK3ESM4SjnIodHQbppUda6QBrlwGP9NmkRYspRVIf+Q/VRDUvhwp0mjhAOyqczbxxm1
pkB6FOyVnE2YuD6bmvCwUU1VLCKkNN24kVkn4a/7LI2nZD5iZWZ7UssXsTUkif2sjg9DptJUZoDZ
yybpQuK52gLM0z0FZXbKbi2plqldEcG3W9U2QcoiWCaTBTa8lqZ7FvpqIuWolboyVPrfWW79ANQ3
p+oG2BQIQxy7pZduSV22MOS4ILMvE+oKUBhrGWZ1rCMm2kp/tbrqCEKha12R6OVaRiuMfAW5RYpz
QwBkj99Y9ar7jJu9rcSPlFBcmErjWJAOkpJpIiqWkwJ9P6eBv6xsd+eXY6Qaw6WwwyLFuyotBbiJ
UwuA9U1QFmROpgpVAfBE9/DblPl5l+ffH+X2wYpt0U2f8kxt9yySOSHQukbXiDeU6/0ge0CCHOcp
KBq996roywQgkGmoXPaKQ9Qtdyb+dYCWlDy6GChYb22vElmIyViTmueS2NLYCb7Jqf7FnV6o6mSL
Sy8gxUDnd3Y45XAkg655UTZER0Gn2NQz7Dg0hW5ecVfwc5S1RVRH2SBTpc33yIpkcTlr585fb4ny
Kx3PUaihZDvufgeJt3FRm5Xi0JuAypsaAv4lyAhPWOZI4gzEkB00K7upDkvLe6gVdgPt15ytN6ox
YQp3kuA6sqjW95/gsAQZaxi4LrLrPTmoh4UB4kr/Yvv4E22CYreaH9rTQiDYJP237lSM7UcnjVxk
IqXZiyvbvH+Zh97m7nAHv3wBYelpALRTw3oCn7w3mSShHOgXoPyQzHoJSMrwbPwQ0xnvq3qBunsK
QQD8W4+bzgxYJ7AU8wqI/iv6+wUMvK4afPMp7WwSkPY5MUN6SR3Ka4/hofpdE/hp7Hap1pErUEQV
62tnSoDH+hoHl0Q4q2c7uiZ46TrJHgpNNxM3jHOXDqQvJSBq+kOlRm4m8q9i+kGwUB778mWbtUVm
lj/P8dkeqcK9qfnG8vtQJRdQwcNzN7cKBEXO76i6b+PpdWrnly6XdQXuecDJFZ3MsdLs2/2i9+xk
hacnpE8uxhm/GsJMBSKqR36q1/wRlJEp6OXnn1YZq4iV0hTRfGhxXUS0thFlsOXoP8zMAOxU+Beh
tM2aii6fv56ry+5RQwfigLr/uf/2mdAo5gOHUjczUEpxE9C8cTMNa4GG0NAZzL1IgkGsILJyh5sl
OV8dhRQHwiKua8enyJtLMdlut3gvSZLtOMR4Iy1yDoWENVh/DMd/lxGxcUFxiEMw3gqI5yWZ6WcJ
Toxr3j0vquFCoCxNQZk/aXEYX2YpbCKKHmq/valwlp+kN4NTyPNq0mguC5h26zXVp+belHLsyLYi
BWytDdW5Ruv4xTrkgtFE6MNAvrEqDGJQA0Z/l5uBVg/X8oVHPtUBMbRMXOScVNZxZYF4YntAlszl
CAiOWoFyOjj9EOpDg92CVz3RDGL5AkWI2lXPd7kb9Jf27d/vSMOcuEGK47pFdiAiaRbnUL+L+vHn
PBPjfeuwenG/q4O3Ja5Z7caDulZCuj4GcYKPapyrm4UC2edf7XJZCA4GgsGRejAWbOFUqVzSXHWg
pTY1zYJ1mPz5ZiEYEedSMdqJyvDlEffEZTZQL38MArJxFmEVtpbJvte71/RPwHVZgu/E7zFxNeA1
F0MISB+hbrtdfJOsBvKXO1FPrBhd17jMgYDLz5eFUXaHolRci8mn4YgvN+aqOVsBV101zDlzDK6M
AzxUsWcYJkXXLfkWVy0kR2cilNvzHYFFZbgth3z/BHwHF5Ar+Ba2F18fhBP838cZw1+tOMPx1VhW
t661Gc4O4OvMjZGJXsGEw2CKgGq+vY9Fq6df5+6UIDsTebAr1FxpStZO5T/V/mmT18Bsyob8155T
H2iD54N02eCETGJSm6b3wr0Eg3oKRAn+kiUHAt1opTyFKlfOeigHS21WPqsF9iypqjeEiqrVUo39
hJY22T/DILk/XuyqKl/FAAkPSMBpC2gRs5q6blQWZk3scW6i240Qqf+DYeClupm8dnQexue0Jpzi
GC+0kM275zQd5V0PHZbynJmUx8oaakxhP42TfAVoZ/doY7x0vCHDrDzwTblkYAki+39ulcbHNX5m
HSZshdeuXjFG0mxvI3lhiTlPzjakpIrE0eW9Rg4xJ5a6Gl1BnkDXKd7lSYokMko667OGBA04fFIw
nMqv3w+4NLttfpz634VVT3QAdk4PIAhY1tWCMWOnyMtyNzhvkUCXzMSa+XrY2AbPOAtTXF2ZBbLw
sku9nkNpg34RdB4dbWMGBVBk84UJqT7bsRFggzsWJ0SseYn2aB83tGmNRSkSV/G5y1VvgGR6gVW0
aqxAMl4G1FVmmk96dYwxEG9UtOyaS3HOMtPqGwux/16BBe1xpT2ARPhwnBw7sfd/L8jWKHjhSwQ7
6Zney5NTdlWjbR6fQejbPfcigJ/PAxjuzAvhsXs7XkRMSuTvLaEM66usSvF1pE//yuGQrEcBKWSp
gTFwiAMYyvnYDzvsrNcMgTaH3pjwYn1jNepoxXNSfGOkcb1G1qAKe2t+OVadPupv+ynoeTOwgv2k
Xz9LsCFI6hhPUerw39GN1n02u1FSoLae7aJ4D0X8n9aYFQFfntXbniq1OVlK6p8w9zDfjcSvVsqe
POPOIE/kisbpYdnp4inUM7UEy9N9MNUBud18bs6kkyE1ngc9QqdJKDtTAUEg0vJPlkG7HlFcOzd2
GUPp78rjl/uOgEqinPqflJJgzxp7sQ2y2S2l4FGfDltQuF6wbhPFh5X/djFQzLprVFlqnxaZCDZu
LqbT/c8YWnifY2BLwMN8rLLD0N0uKvhnj0XSEYJ39+OUt0yt3wLVGo22zyQ66KJ7v6XqFDs3WELK
H1+Y7sbUA/O4xueh8+39ntS/VEcgkGOyU0NJ3+qVfzF6/LJdF/XiawGMYpCkkJ0zTUCuoy6nU6RM
+EQZBQTeWacYpgvcpBOQy2EJ/9tbjyaSX9OjyfNFCJZ5nZbCYmdBp5ImVJmfe4SbaaDZOkj6ZFcJ
WblYZIAy+aLKa4iKtK6PKvt5gbAa3N8E87EF+M4eVXpDK9WrV8+WTOASgWnPAt5KRr1FuKXxgbtI
FlFBmwZQgtGn5mQuqcMexGgTMExxWhuXqFHZDeBOMeWQdLgWq7jlBmXDAdamwGnS5SYy78M0kY0B
pp82xWmpVmC4UMnpfx1GcU809cG6PelfMb0Kvu5JWzGY1ZSOpR0MdY/KTvMfW4n0ZClLVB4/PEGW
5XmuHXjWJhP2WLWucM/SOtQoXqIsIHno6SxXaWE4/nkzWECO4caiR/DklCNhFPtHCWWocmPdThoy
HZvc8N7NK42NjJpoiTDcAK9GguDsgL2oUv9hz4w80E5M2KxmRewgv/6j5sBXKbQ9T2AnVjZEcffn
pdeTUkYGstL5ztYnpwDhc2YOSJliVaoGSGMj90l+ckIdMfKcTGUxvNAkqaRi9CFJIFw0MXjkHeEB
89ukTG+tBhZv3R+dCubReYkQGlCpd5yFohvRi4w57DNqmsEYGIokhEcJEtxTbQs90gpUE72wSmiX
L2mPOykvj8ZY/ruCNwuXgcERrHBUThSuW+ePy95h48PgJ+RZL2111M1+2ar9pw+9MjTxd56duz6U
kQ5Q3lfBZrIh4EkVGlN4RFR94km+DpFLFCupQJklF3VfI/NgXhCdcPMZT0ZgfxoJJLNLkLz76YUZ
SJ/g0gXuLMjLfBSEOyNSK1uc9fbfDHbIwIcDukI1S2udkFv19G8LxvjPTqmM78b2x2Us1Wm8Ohu6
ugjfeUgUIPUz8O2pATB1FWpl9ij1L6/95Mdx9Tvfy+kr+mbrPU86CPfkczv0LEd8J0JWDcYYGKYN
OoXVgZYyUUKDPunX/fhRKsYcoSSCqbRmuRdDDTXJZq4lVYOlDSm8Dw88o3F/iaMaqkX184PHmNjT
TDZGPnJLnkjAneSm9JaGLPBQ16akzXtm+byOcgaVwIrHUUpPhlm779iYc2rq9FZHmhZJc79yf4g0
DZbX5kRmydbtvGiajGeN6NqH47qA8spNdCUWZGeIqU27NK3y8EuhDC2eFUvHOO6H7Zesr64eIMlr
8AxlW+Fwb9U/rmFrdsQj04qHnpDd3sjxx9k7/VhZt7YR2UkZL0bYnxZCySZ1pFyGYBnL7l4Ns5/B
QKz2siDkjl886wEsxy8A2HsLu8zJscAuTjkA4kORkfIrDyRmQxjj+6DsU2T5lIdkC9+5et+z94t4
VQho01ZNTnZDN3ZwRf4hCLOeB3lFdZttbG7WvCGdy3vBctndOG9ycNIfx19ESOh96y/zGETZ2O3j
hovYTzEyuNQDo3IakTaf2TvFSvEzuY/nVCuwCjYFaip7MWsl8uWv9wEoA/42xE8NpES/08P4vj8t
sE1lYWhlFqbLSd0ixACfD000OhrwNe5SjmF/5B7Ig6PZZe+cqtTvC8OHYM4g+FB9Wcd0iA/xMCZO
CQ36t9WDalu7C598S/o7xRNk8DYgwAkcqGEFfd20nfuEeAHnHJ4+etpUol0zQsARJgFB12Ghcb91
29HCwtwQbQr4M7NolOzblvp+LLMm4HUtV+6DUsTWrVERRH+g0dxVM95fTjPMvEAlmLgafymBacl1
NPAp/ITzcsM4N2etVoPWlfAb5EeYtRb3DU6hr/NoZEPeVkU8t958/9vfBLe1wEiuhBrMsqgctJw8
jOEoz+NLhXmXDJJkW4NZPoeJqBDBYhykSWHAYuuxRkQ+/ADKdzJgLzjXcR+8HLA0RDbrVVoSne98
JiCXPJL6WA3kkBWIRMak7kFcXXOh3Tw9BpLFKA7sT53s8RXCkB7btW2yLlD83NmheGfgDcAccKzk
hSrgDqnj1+/TTjJBYFnda92wKxoKTG/HhFcgJUNAiElcSdYqoK7/hP6biXyP6+jwAxQ9A1GrNYEl
GytcwwV3KtiISoIQqrBlv6I68kYFYVL99oIapnRxL3UwBqr0my2Cgxvah/bRZyZRQNMSqhwdCRIP
v3usYpQuvsaM51P/RLBsaZyWd1TVroMY02oZzj1DLOxWnboc9KBdlSFB0w8UFI206w4tdb1v7fQo
zlkACQWOjzm4CvemUziGkAiPi9pwvSdEg5MAQ+MDdFzlxdIUIzY0YqKge3lE8q3qFwPRhq068q+w
bb9jZqkQevhgN29WDfq3U1NPeY8Vb0jmOy4ysbaeKSWZwmEtbQh7HQjCedKQtpjvJni82EmyjYug
/YG1Q9xnZxsStdQ0zUxv5F4rf0iRfI3Nc8a59MXy7koIDucu6Jw0LYSba4hgBdk0QFm0pbaJY0wR
DHqeh7jHNkonsXLQHeF9QXYtHXhcnxuT0NjS4bMCBkWocqUD7bcTaJLGjNuRHefvilrLm1pPcziL
07f5EbGM1OD/KmS9UuGGy2XVLa6LdmmMgB+/GeVtyCZEfjiT5O1gd2i6i/wAt2+4dgyFVpo0Uivb
xKpQysfwKSfebh8AT1/HqHfynup0ulG7PpuwCRI6eryLedWmyfZwm+8zAycdL60I7KY/bcQiFUny
fn/C8ZTDC8porcHQd+19QIBlGekhehAMg7IXj0CKwdOZYTGhhQqFvDpTXbJWb2h4nZGWq9x3qczp
PUjOl8dSgDzZOk/s/x0KHdFazXXqZ114PRTd41mdXpDE4cWShfa9pOgqOeBwLv5p6K1NZxRIbDeB
jmfdAgWZ1hGznL16SsvapIfg0tTeXlXdPp6ceA2pdmz74gRRL4n/WSFrYhEDfXFKwGw7WFT9/hEO
nuvJSUmwDk4vZEIOmrO+u4Tom8UMU3YqMSyhQaq3CAjTc2gAd+vGMSQ1z9HJkHiQ9P9tjkSJvnk7
u64/p4DiQL5WD3pdXj7Fumlj1W13WAmT+Q181xeg2KJfuumYjqGVgnWS4CgxENFRo3HYzLrXFSUX
WgFNAHuyEijf++crJq71Yiqnn0+/MZzZSw0yyuV8Ub6JWPsW1YuB8msoRItSprEMwL8YbYEa/XCq
oIEkgJ2/DtZfp4YS5DytLSVqgvyQY7vNQrn6HPTiOYMV9d2U1b0kDV8RDOESdiRQFNYzfxNDrv+1
poHvWR7nSHC5adslp6O05uJ24nQ21R9To8wJ8JO1JXp0mSicSU6q+nYmNh3tm7U8Iggdki3nWQZi
H1zqQWwINE5fhkzJQ+rsbHoPSaBd9jWOhSe13lnrYTONXKxNoOHrkSH6kcYZnEuLhsjU6qATLxbh
L0lW1ACumuuD2d8Ooqnf84vbazhm0QbigwYNUZk9xWrFxG8cH9N165L6RetHwuCeffsMt+9Tm2ge
T+voPje3Y+ufumbN59swc2EtM12T1vyXkphiz5lT/NR9DcvDQ06+1kHGeyCbZ1eAbmB40jWrGEuz
g7FPlABAnWkqythVBKNVhRBCBEgnwsvARmZdDgAsVNaNt3xyGXAx8JUT+i6yYPb9f1uNNAFqUVTB
DED2NcII/T+zDyMGyejJueMyzsrXkjI/SH3TqVWMhQNVZk7Cv8QAVzv6S94cpy5Oehl1QHUNrjwh
kTEVQcEMydu4CBgUrj3/1T1LGixDiH6D4ttyUMuCdYs2z+5vNZWKCThXW+1+blPA4n8wNpHJp5sZ
+iSQbX5H8LD9lxtW01KqyG2KxWy7litI/HC4rZebL4Fix7wPpqATzhenddVYgBSVEVQr1GuHf7AX
7nc5pfKgTpozMSBOfasZuD0pKbCHJ4te44LHxOF+oeusJQzqcS3QYeCdaUEYqxNStvCvA4YF3/0w
sfwG4zdfIFsKL9MrhM/iTwAgv+7T/Tjagai809NqeWHvCyw9ihzZI+FshKkkc46LyauHfWs9vxGm
Ro/e9ID2QUcFMlgTaSEeif6Y5Mcdd9HmT7mVoqntGOE1nMRQ8fj+V5xW9qBuUWQrHfmPhwxSi9GF
1NWboWGnlguP7n147BxZC8Gv/BdXCuzGawh6/VgW1c2RS2dIxej7lrwEevXOcBSqJ887a9s7YQhT
sePF4TZEGkaWLc/YOM93rX14jNaH8zPJwm3TrNOTuVfSLSHLuhTl19iAANwIgA3naJajyNFgcBX6
0SqKUqyIJ6oBJ1oX4vWqUmjN3JkrQBLzaROp/WuDyTDWLm6aPdcBNGITRJgh8zv0fktAbAkKZYym
XpKEcmYhHsxSncfMKjNDYwKoKUuETnqzdEm5SYei1r0MFKAq3ghOghHScDDS0f4vSJx1sQlB3Fds
USf51iTS9CG9hbu5+P8kqDsh6/nridI87HdNt9GFQvZvyzfIEMqlui8+pAZsdGG4J5slxcSn9zex
WPQKNcwGNt/ENrl6vVfYFKCWm8EZcGBrLAGOrVjx1xSI59cU/kkcfstd9qGCdha9HA6eufzkYg+r
XMa/0/2izLbHclPHCB6lk8eAzU0sKnYxqSQDCooKNsV2s2+oadrs4tx9iAkWo7Fl4cQnhq80yVs5
h/K/M7cHXQlo3hTgnYLz0xWR9ktqHrTWyUAckZzwfm1VCuts5WTJ5KEhprZ/d0CPI+npWxA7PNRw
Ybt3vGmHEu9+vNENnxvIq336QZEMGiuDhnoWQXxntIo4GxqGgJGBr0y0W5tSxOvwFSFPu0+5QWLe
WRmmVqGCjjj+jl9m1gq+gASaYRWYm36NyFI7RCqDHk9bNpN3IY3dpe/uLnTbys7pM7f/eYU79z1R
L4zxsPjDEsD2v6u7Fa+RA3qWb0EgZgCmUhx0x1Q4f4u71HJygIWlJSUqU+jAYx8fpVjadk5NV5FF
YYnzpJMZLLojASIAOr7rMv2Clif9MtvzVpMBhuEoHjJ/V/ESkGZqCYfcc+n2X7F9RKzNFkbbrMeP
ssekjZCl5GbPCCP3AK/CyO+1MA9U1OADVH7yq9DFaFGXfOsXdFnlcoaSwport9NLn9SuJnZbJg83
/chJQ88WVT9aCF19IUB81FPkB/yX2PL+9cRQ7tk4tUfvOn+QpgPb2xiP4qeRQmSH4GvWOSIroXXg
rqpBYim6GaSqIg/fYRlHnQW7K6h1D3lrS7hAqmXDNDpu3wlccz8Bo85nCDEeGAklUGH+UuffKVam
fVCCnm4SZWabnlCtk9QpggLHrFRsRXK+AVqx3v5ppbns7CEqmnBzphTDAgejVF9aTBOWebllEn0R
WD7oi3fNvwZfZeff6uwJeuBitDXyrsXSxFpuCxKAddqnwGnJY9QsUrurG30PmnWgd17K2i/LUwjq
Gcz/ZvapvH9n0GygVdnHaoMrHnW1g63mbONixatzB3m/Df0hWTrII0pReWHvrph+BQDefwcPClwE
zEBBLLaArJYDfWmyqbsEWf0jXJ9r5yut/5wgCsTMUoC3c+AeeEgR3r1FuzCeq4VDegwLw2mx0Hrb
/kx6c4HYHp1PCrYvnfySlmxN9Vwq7UvZJj4FWwkMx7KQyM2ijauW+KX5J+xNCiohojf8JXRY9NNX
KbgCfHeKDjcTXQ8dcu/8hZSpQlyb8BWFJFhFGehmO1Veb3t0kGw9FSfGrMpqXSg/+6tpB+yUBLTz
HTVIbbWpr824bBCo8dB65axsny3+sLptU+wcvCEzuh5RbFZQdCRUpKs6UHVwcnyOe3fLMaBf6vX3
+so+iWiREH0iqHU/lbasCOHBRvyO5Q5nlZbTqG6lg9ZNzFX0vU7QpKeBUBi/9ccJhN1B7lFMb9wD
ngPfJz+ooe+TLrcxjyUAT45RumvR2ePt/dw5QpZOgtVgkv6dWF3gbtc+DQm/cSzqApotAW9ESz4S
l3ynQsGP3dD1dfG74k6U6ZbBj7gojnytVnHTyD5YaHeVmfh9ocPWQd7N3aqY0srqHgO2+INx4cBh
qfSQik9ZrvxRhH1fGBhRZcPG8XaKvAoLg7vrTc7WdtY8ZepHA4LldFm+GH1J1QS/YWnpLX4oUJI6
33ca2eMjifDJD7LWzTMSUB3vIGbib1cCNoa/so0uMm8jleq6HnxeBJh4pfkYletEonbbR4AzosqX
P32ufATzzQX1Pl0JV3aijppjEG2mm3lq81pVgIhoz5ULaw0lRxAuS1bzamDPa71wHSu8eyqkJhau
7wUs085AamPZGMPzKgzhK1zf2JPh2248hyXdHcRWKk6e/INy3ZrrvlezatO+rglamMeBHEu3B4xQ
Yzk/Qa2arkP1IGMUwJdPlnFsw1YxGUGW1FTD/S/uDedC7Wc13gF4Imlvup2kmPGa4CZmevUVxMXA
uahVetYCA9XyBvr1b2fHx+57u2O3kWGrLBRfFTtIZgG9OlpyAFZW5p99aOS56zt/dbGpS7UDpVSC
cKKf3cLSHcaqw+bJTw8cha5kaI1M7jK8AwsX66b4AJEGruh9NiuNhWvvIftnZUFy2+saPf+szCh+
HKz3esLIvocNePCklym5vw36eqiB90zU/4cZgXUbE+2ioOCyHaKzaQ5AFnnpwgW1VrQ9kB18n8z1
+iJF5iR700RuVyh3p6mCCbYYekT73DD5DXxlvUm83ZMbFUKFJL38fGMQ61gBK2dN9PZQ+Jyfn6hZ
40sXy9uzho1B0+u6nHAEeFvqkf/Q62COllzlqYqPeh6p6Z4nK04E6wjCVHgE8kTQL1KjeFJbB49n
/QrxJ5MUKsqH4DhfxUGxm8OI2/HPhPjqwcA1nMaO5P/7HYQlt0w7dU9TGjEYEmt2oO2/YRrqNsj0
6LhAiYARfMTVREtD+tAQEJe1Gjgu8UBo7M/PaBAJc1tgYRH1EZ3jSKCIe6GK+Id7kzBsQZtI8VuB
Z5kzz9V5UCZuF7JuG+F9xNGugDmb+PdzkiqgHHyonwTb0SQoqklsTCtY9XfY3HcxDtVbfvUFNjyO
8URZ0hGzteWh/pEeCMFrhW4aj8IEFHmbmMkzS53d3y6cLROFYVDo4jeZE/qKtyy3gfrfKwSyXC5M
tebnnv4dxskQQyFNPMQFyBN4WlKDC7C6IxJdW99ZCRc3PgyJeo0dWAdZVJG2+HgR9CarNwz5hg3D
DC49HZ0sJVbUhnxAMzurgUzLFy3cG1yB96SOSroeBL53xSflpbFAHJzKFgNSa4ZF35QuSobr+VKQ
/clAWAwv8fjdQN90CaqbsaETBLXsjNXrC6IxKpLYwY5botIyZaNu6kAbscfUUBPoqsHwrfsXo9US
1oUf0OSEFby2rWLUdzNOQZLM+QL+nfJ3qVBTOGGpeoZNJpLJVzX8VmRRvT0lT0DDgoQtG9/60VXF
iwqMpzwGLDzWBImgI/1vJljZF0ky5jgrHTzndqYyyz+W9mfwwChK+xOovkNIIRCF3MQGRTc27nrq
4vVrvLPnU0ZGrdP/QrfhiOtMj5ywQrMBFKctW+AbU7HzdhAHwQx1GDSpJASakf4YWUk2u9K3Qa0U
SvxXP1a9GHDNSJ5UXo2y7WaCKEJKeGqezaFn2QV69guJEZ4sUgPpQ+wSmD1fyfQvaHx/f+Xaap6U
RiQX6lDWpRQdG6n+S5X6bFWLS3+aVUrW+E+QOK8imzfkZsC5I+JGeho4ktgeKDaA6rPpI7fMZ8qg
KgHt9u2lck89J/t1a4Zpi108GjcEiFQ13afSzwTEFnoPZ/CNVoS0NEHbywM9m//3k6khznzqLDr7
RNPxwZf8oYvRPJzpde1Ax0+2riT9XhKiv0fXfVzpYACxf05sUtCHZr+JH691vk1at08wuV7JRoQe
3ztILr76nOfWIPuq7gBKTS35cl0oLLqDbTHP8Tvzxn5Mv54twyq+h5LlcNbNbVDrbyLVld9YNMnN
Msfn/O/+LDfjaLYTxqadgWZaWt4yVc8sFGcO2DvQmAFUw6RGqCu9q1C01d1qmGnmmw9K0g/nOKJh
GelEGqSrKqKzKJ0OIWhI4y1TfV9eWm6ssU2eL6k6ApXO4chjJDW+RPng7g3BsJNKhapYVgAnFr39
5Ojd6WuXGdUupD7NM9qb8LElMNhJ9k4DNK1s9RtnNMm/HZoWAmKVySaa87zb2ToR1I+v/9wO1ln5
qt0A525pmTqTRvo+9sm8B2flxszgki7S4yLdSCsRxV8RBAAK+x4wS2wTMV6F91pYtZmL9pYqRlNg
r0849iT/X0+TDbI4x+zTnqoxD9VcE2fedYqAQH0OOIFtYFtNxPzm1VGCTNHLdm0Rbry9TmQ0K1xX
ZxtJSUWhuivE+bibXzhLNH5X6NwqVr3bvEuYua+amWEt++6tcSOKcm0bzAfLtQWyrcL13odTrATy
vzZdrY0c2IEybg4SHdFEHXcMrBRS9V8hSUtCopuI+gEqVwYs/knwT2BRopMAmvQrTM/fAZk2mW/C
NPGC1kSagfg5KFHJEBvxruk2eZsOKKY1Z3ZjEUj3BDfEGIfq+0zVF7/30leqN/IDL9wwAIxCwKuF
pVgr6y+yXJ15pstEhIcqONeTU+Spjd4BFKKZ00FytCIQ27i4TnT8D0ENuxw8UQ9/NX+quN/vng0+
g5IdTXRb8OhUdIElszVxhA4rkI+8EWsiY6CBAqle3v3At7LO6/3UDbpf+RhNpt7DwEj6sBGA/5uA
kbjSbEzaRwc6jIE5a0ZcyZrRGS11lzIuK4glyIWZfityTmV1my5OFkcgrRRr2aeYrFByZf+j1LI8
xZJN+kqAsvPUtrn2p4HalyFXIIa+Dwc9qh/5Ww4bjFklI5GK0lzuLEzg04dBsyz/ZeEhe4W1HzCP
OTiPmIL4M2ndGgAl9vw/DjuRb2B0wRMXQFO2jVZQ3o/SpKt2D7a171MDQ4oscLjb/5IbFltFvTmG
fVXhQFuy+rmi12CvsJqBRPNTeMA6iaI+cGDVNcbZxUUFDHpzNI7wmuoXB9yEdCuLmDYntWgRuQyX
NhqY2Fg0vM6My8AMqn3HLVSBe6+gxiFZ1aYfb+1wIer5TU2sxfJVjvfDxDYosP2/PK4DcKjgBHBc
WpOK5zKYvkgjnhdUfyUGpKsBVwJ0xO823GGCRVhdh+l4VMwqxVYiIpr9nsWaB3sKZNvoh2uz5C3X
N7cFkrK7sNzsXcDfLL54HNBryer307dIKYFiOc0w7JL76qxQKvfJ3+Jl23J9DQD9d7yZ+6naGbA6
gKMNYFV9nYH6mLZjycMvdbcjrYINJYxxCsZfVvkCLcjlZi1+vtrQ05orO47x8zuxqc7436qQwl5Q
ntXiio/G+TCTZFHJWecNj3MzG38lXXQoQ75vFxUS+eY552M/xpMsUQCERxRX9OTBoKvykGSp5x53
ylzUCOPwR7kc5dHZF6uqZFYSzv4FDE7cNpCrWYHXX5Sa0CvCU1ZBTLsGUdrYXLVV+/yLUlPXZe8l
FgXUfWrf6CRwwc9rBmf83t/tzKKQvdVPdPHi6TLwMFaUbJjC5PFQVq0j8KxdoPT/beq8h1039IKN
MKJKtHEj7rTWDk9UjFUSlYTTjPOnAe0U6171X8ZFYEYP9ycg8/miGHJOfTCbY3j7Q4w2fz8DXz8v
Mq1Kp30pRhKEblkMom6NY0nAlyu+rnDlXrutiQXC6MYeaBQXD/p63vK5UdgzsNOIT5Ft4MQyDZuX
EmJ+YX1H8kaOj7WBnQI/00AD/0/HJ2P+Ws92RNL0DyTQ3jRly6gQqkJLqWhqKwq6x+eVWlWAooAa
mRdhXhqw4IzN1LNHqwTBzuDk8C1J/rOFw7PHPdApsFs0fT3cEaYi49H7AXT+AzgyUfRyiWV+WgZO
CJZnUr/2UU9/Qejevn4ZBDYdp9e0FEJ9q2eiH6iXGfSmCioJ33RSZlBP/pHrvyoWCn+GPi1yoAZf
cKAmgtWD3fhPvxFX+dGEaFExO3tPYJmOS69oVdJyS76XgVVKrc9qZbhuM1TvTc927476GU8a6dQl
LBfb9qWi+8q/T5kqubawuqt+exNdfpa8SVw92fkPHIQv1MEXUUIV/Gn1BJSKwKLf835eB86s4hgZ
EodwIkwjTDPsyAkue8b/edoocWbOlDrwNxHSRhn7M9J79I8nlMFayXfAqcjF3p86gvEX1aXq9RJc
6o01IaU+Jd+y5JN/VEsZFkekemUlhVIC7KV3eqpzmclVSGpoRrAUDtFUsRIEJsp6Fecy8ZAf6MLw
7eTv9Y/uP7SxedtwgkDlPYsgrfPecoiHDGcbOZ6/a07VG4G7U8LCLJvHA1Z7fFBF6JAJujxl8Hq2
+3pEbTOgP+N+S0ok44dE8awp53MMxwCwAUwqkW255/M6pHT029qUcXw+/J/MQ5yNpxmNSB6Fk9tY
Bn/0gHDeSTcFO3DZxc8/mEb6l3WSa7fWXY2GE25XWEqjy3ze2CmxL0l8E+1C54c0iVmiOTh0tfvj
xlr6Nv7h37TgiE9jiq5nCevFBYptsaDfAn5npsXXLhjcMmoSmpHcG0Rg1bOhpb/NRL6FEQqk2fAo
Ry6za2zs7YBjmMuQi8DNAlckc7Y129kqpVkkJBIfWx53ZpgFFI4PwCkYAx5xXoT3PpcZAYH+nhNX
QnzPCB75ToEPFpUf2VwYPhvYOY37j0CWccfKi630KYiyfA9wOI25FzOGu4hIIY4jkl707kjzprN2
nV2N6kgV73GIrEkz5lAiP75m1fdb6qGqt6P6+xVWUjnoZUxww1S9kQdSPZR5qbQMiY1iX179wbdH
h/GUMrToBqZzoukEEtMLiiTw2/JTiDb3eHssiqfL6LUEiweZW1LrxENk5ML3vd6R9zsqzl1TLaV9
y5XLhY7VYzxoFOqgw8QjKKYPFWeUqoYxFG28oI65vtkdswJHbZFAH6KLRFRnFklJjp0n+aaBsEsS
d+runHtfhGf+pEdf+Atikr/UcxwN1goDE2qlWOXsML+AwhFrydewwXZFNc6zL4Y9JYWx0er4RB1Z
4gIOaomkl/XGoY1B3Yqgz4S9JFq7A41oslz1XHufBTI7NjG9iMvo+QFv9uYYvGaw/p4Jp2RVgjOK
oPwPrHVQ4cTtih+8CV9in7pwkleC3NoXyJVvNmFMF/5a2uT+0dChC3+8+OSaLzmeSD10xPipmkOU
Afrtpi0sVjdwwek4lC+fEZDLJEddJKUaRxBmhtAXoNFGraa0L+u2zTmUMsymhabIbWmgAFdSTvOs
EEjlLZxVs2pNDH8JIiWHRV/xViIdJR9/dRg5kBK9oH0MHSsFa8dqihTJou2amfHk5te0X0KSp4YI
/zsraGjRokkVckgc1oEjxCNyK1JQeHMCYNtY+Z68twUZFlABEWyPNijUl9YuAh1TZ3GPFhx7pnOY
i2zIaTxxW4Wv3VrL32AgK1Zt2Iv6nrvwe+bj2TbQaVsyjw8BYYDU3HJBYDTOPMwHYLt3PYzX2gh9
EFv3kWw6JS/EuYDXfv652lj39Sa7FvxTZrVk0lbx1xnFYDoGjAQXnOAh2qclTG5da6sNGxpst8Nn
ziZwXQ0jsfSq0PUdMhkZNkAsxj4cmpepK8aQqylzU6LiEYdaKV/6WPxTeHfjyEUYyQVjF99Jl7Tj
ji5KKMdxkNohtaNW7JWdDgIkvRwlV55og0CIQir3fGn/H/CKnYKKmfK0XN/Dop3YfPyl7Lx4oFUF
M9htf1gT5J2WqowDsFErWi9LrcUkKzJD3rr+O1CM3S2G+ouqXeubKjqBu3m26OZGQMYfPvO4AK66
fAc4XEgqQbfWTy1uH94ncz+RFp3+AfJUNHze05sUJixUi/DfSxaRPpxjGa4ipzARiwAJlvN7KlDV
KiWhXHY9numd37vQSdubFyd9ZXT5HPyjz6yi41P6V9hVLMsWFOgsetIXVus3Np8UdfiAov43lCw8
bu3oIMhiqufaj7uTnGoPbCqzEwhC+UOeGZRnJlqbZEc1Tx35sC818o60QfP1qwTkv61ARkoD8J3h
1ImSKLSPt6Bshgj6EswK+JG5N5+UaBbwv3J3yz/TnFgP027Bz3OaItqvOX5d+OtIxtaUwJUafCpp
VQMnWvQd3ZrvcU5b8nwdSyygHcGnAWkAUdMZd9dODrzWfkY8tipgMHnBCUAiMBkpSxLoUJcfNqCK
vJyU2SukdZCXkXHA7wHGCq+WnbQcbDOmMhVTVoPdwgCPcDI64AxyblCQzslM0IYDswlkkZwZ2kXM
ieZiyIJOuX2LxZSjizMxbPpN7MtICcgytKexrfI+WWuDvisn4KUk09pHc3ys1DPH/PnZUOtYXy5g
uWRyEacs4J+9lNHTvfQarOfCa4m2FSmyJfBbx/WmQvxG6GaoVeL4cskGaD97gKyhSsZHnZbADLBp
xFy9N0X4pe5+/NJl951Q/WMq76sasV7eX2yxuu8KeSuXxwfStZAc9gXP7cKXhhZDonoRDgeqf6Wh
TdeZgMZbMo9vYDOVwFzJ6O9H/ikbng0GKOTsUcZ3pAbyR09aWYcO/vH97Df8H1rYgKju2F33M1jC
qzFLh4DF7J94UzVQU5PUgwDVY1tXJzagdv0tGcAecEIApBS1D9sSUbAj0AumN7OEO9q6/A7rLjCD
kk+wc8r6VMLCTnTV3kkKftugpgB45vqMSG3Un+TfKUf86kmra2yvYkd8SpUOC3k/QmeiMXQ2ZEoy
c1tzl+LAwJmj/nZLbQH1A4vXBRpoBXnQFEyeH2shGiljLK18JjSFMgx31KJYXQ0uA7WjKRJlJnnP
EUD4ss1FZ+cOeV+YL2KoNevEs6i6rryBT2LcYWR3is3rZD4EzChg7KBcK9oJ4OlnVEtj+go/NeO3
dJWF5LQqUVQeZMZ/Wu9XiTd4t1DsH5zKk/GbV2MBiRCB0//dXNCo1W2D7k+oQSTjfJmI4UPfbIEF
o6eRzuvWvrUYVq11ZO8U0Bx8aO8KH8jLb8VWhqYQkCrS+dgvoJz/yZ2fzq9XXU4h1/Bpi8KYDuvr
JZMifi1X2tEnNfG2vkuxRA3DG7SA8jDFhZ9tW4lIIXwJrHDVjBL/gicJKzhemjEDYnyK9PaZoseR
hinuuL80iN4DGp/qWj9n8doaZkL3ssy8LyBOHfaEapXJnz6uqloIfiY8l/pw2LrUeaURHDgUKGEp
cJCXA5Jr46Z+nDqBcmFh7AOQqeiGGnkHpKju/eLZFfU4Jd9zY/W9b1lcYGd3QuVaDrpBWMQQYrlw
4wU8BIpLbImDklHNcJuxAriQucC0cdnbQGjqrHEO7T/AfO19gu4Z5kJInCLxbjH9+TOROcd3jkdE
HvBrl9n8wBZzaUcpknsGvndrvL6VcA1hz3rf3vaQV58KOr8Q2Gzmx1r+xVPJ88LzOLRnS4WIcWWv
AzqgHZbIbOmTi1sHIQnRDP/SOGE9llIDC+aQ6QxA3FctfVInvQGsSgeMbCyGdXS8TQrewMSv/8eI
6e348a/cvkfi7sYMdZoEGJ799/hg2jepG3REF6WhD33hjIr28Hws4ZtTaRIc6RJWy/ZJOstoff5q
fYchU0xW7WLYAgYdOuit6NdfS1xKC/V8spvpLouH8Qs/WtUe+T4zWyXpTNnOlSFiZfwO9GkjQ9ia
setBu20nyOuwm3WTjTkH0CXIGbmADqhs9LQMzLZBIWKxbmyuG+cXldk1F02WCEyPMAIvOH91RMv+
PxxexRlGlzBvGgGYhVMhgwum13UiLSPT4h7oVGZYXoS6J+NBRR8kpeCZIZNz+pBtU7rg+tqzdayf
uZYIl/YgvKOkLOVQsOJzclwiJQ+7bOxdNWEYQDMRB0sNcB7TsukEdwVU13s75w0yiNHd9yQ0dlsS
GzJLDFBdGBOJe3Qog1NG+0yuuqxHmkiTKPL36xSYbRLKSayUCw5KviK45GbhEWGziNs8nNX6/7/D
OKmW3Xjo3Be6Nv3LYJtIMZui8FIMCnayK02hOTc/76uaDy8fjZnXLXr04/uBtI05LDfH4oqrDyOS
CiNvRP7pl60C5rnBBrRfGtliQuocZiYcgm+IHfADSz8R2rkA0gJnTziH7nwZO/UolmWwv1Q6WERQ
zx3SadAKAgDYF8AkrSAqo7H6JtAcvQ9yxw1I9/8+bUDqr9KAjlIXBu7udGltLcYK2z7V4wsqSX4h
g96Oxv3LaCEcQawJTzi45HrB0iCZxuMzUHfPqOw12FIJilkB9181eZVhRCWS9P8/QhB3S1S9tVIf
eX64VjX1i+0lUJGip0tnuMZyMe0uJmLGOw1on2Ns/pAQ6LDR31ZZzWZl/3bgBSZaydt+u8WSsIdQ
+LOY/fUCq7di1n4OZvap/zOLboFYgWDuV+wXbpSTqPFYpcjEmZcMSWO0sCq33yBd7yVdnGmSrkKs
owOxPrjdkA5Tt7m17zwkyB43ZhxhIVZiHW//czaJfPALrUK30HP71k+mdvLmT+za+idcyglfVcjJ
QCBHsSlKqyy2SuE/EL+gVPTanp4koKGkcuFl7qsRkVgqQrr+EoR9kiDZQX78Kk7Zdj13tIFdNBSi
AZ3hdOLUI/BZow7iCvmSWQ2NA+CixYdqpSBB/nw1Os2RN05j2jX1pCzex3PIqsdKAnKiAKfzFfY9
1FtC4VH7mAvB7PD6McedjLz8csC4u2yYwnv2eWFCOLN9P9bILjVx9ybjC4l8mqS3G/toc/tHwF0K
0W05y2PnZrce8tD+XGUFZH7AaN02GctczK+oI2EQLBGfVLh+pfnxYf9BW+iEPraWzNmCER91Cw95
oLP/PUwvSXH7B0p4k5rfUKy1N0249l8tB4GdqHwBclR5fbhTjBGC2a/Gg8D6pUBP024TC/KlYUd0
cniPnnamr4vqfwXd3X6NWcE9MqFN796lkKNZXAnArGOEWMoamxTd49l/uNLVIF/N9j+skAS547Mp
KKlgfS6uhuHAhVe35yEtIMiuCUtTFys+WlmneHMnxJharPogXwA1r/+oZPZso6FQUfYIL/kjXV0q
87YCgrW1MjmiypFVnXx3w2pEufPC6dIxEnjbUd2YHD9ehWS9KpJm7KyGNVnEgfmzb73cAUP9C+Q6
1JEXF9GhP6WHOTTLhqlTLg5n2q2+U0oGqBdCIYcgWN5cK410ggFWlGrpyS8mgkDoewbd2RGGdGvQ
U4lFA77x8oa1Id2FJq29ms/SYRueyiVG9FfLVDLpawx/HacoIAf643bkLnEugTF5fQ3yU3xpN2nT
Us73vfM1zOk5bZuLr0ZQ2sYqlWuJ6U1XdQ0b+Zz2fuwaq59ha98tgZcPGJHJqcucA1YO/mbNbo94
vxGjhOBx3a2Dh+8z9V8qh0JUn8PXOxVx17iljj5pNTn9WA3CucyT45nz7ZQEyXB2R8ZHEsZXU+k2
tVO3EHg2Yqh2oCZPpJuU4fQIwtEb0Q8fNhoN0sjdiY7Q+RPIJJZqIbS867c0R7j0/Cpiq0mbGgpm
vOAThu7lUymFyZOkn5lQ1UGrEDQtlGTUXSZ1ut/ApeK1tR4oMBExFvGQhAfzDtHBEt5fHNVbrGOf
7YZmHR1qrgAs9KPJ0nu9cQtHRxCAdAhvw5rrKx+WXrn8/JtkU1rFS8Xw3nrcG4i6II6dgZYYCIeC
3Abudb6Gtcrv98EkKAIeeDAGDatbkRFVwSut7JvuSvx3vj3kkb7idjQtUEqFMeFbtS/yMjowHG06
JnQ1m9Hh+tlr+dLyRdR0Du8qeWaw4Q7cvleScKKRaxhusLU8aJfofGL3yn6X3YJDf1VSQSc9DtXx
87LS75pcC1vVI0MEdJNq9vqXh1Ky4LW3R2epZOq7zJO5ktHUEg0UP8Ho6rn+x/Z4pHkF2Bzj25fu
28zcnEM1f4nuMVh1yUkwphzFxtmwPyq9df6gWB1r6pvKyWqzRTzp4u1pE5yghedGPKCtBPhOoZXU
rguViJhPAy9asdraD+S8SYePuHyxywWfkji6UV7CJTpd1RnBcjxg3836V4AklglhekPQOCirRBb6
TgwtXLNWpuV6Bh0cz/XSHQ6vQEh3+ryKqjndsxK+tqo0/S5se7+fzGsExU5cWBuc/TwXKBl1XfAR
ZxlhejaZeoklQB7H7Bn9IbfTBakDqwbfCPR+y3mrRAM6VnzgdUbwk7VDN2tVDIdwz4uJCysIpzYe
RnUNNGrXxVxicry7OTs+vsxMet76sgsXsK3p6AnlfEyAAjpS8pEUTP0TFeHllC9SVJbJ7LNGITfN
VlmWMlVOEa+sTiXpO58GshxMyC4QxTPiD+6P3GGVgrHcemSG7gLj1huVg4gRSq51M/xCmUowpcR4
3Ntd7U/OJOnYtphhupw4RJ8xqsf4avRLB+PKfw29Xw8KPrKExwjC1You5fmNayhChOxOaT1ubbmA
3wlWJqkbGpUQkONcW6pqI4+EczE1anvpYhDOt4Vf4JUFM4+jwi8TdvJEfJ4+Af7qJsQgnbOVRehu
HcuJRrhBmaJGbx4BYMAJXg/LmeJob1Joll0Y+8XowBRvHs0WcCHD0DKXju90NPRXtaVie2250LqP
SV7qNv/Zq4o2rm919WNDa21p1fPA2+QMVg+CIYXsXeK2O6W0nx7bSuIgGiIYLxWxji04+MmO135X
DWnewYnaCT9ttPHlD1DEJ0oFtiKkArbt9CJNOO81TLf7nhubDNkoLCZUC0ynFbWSQlPO2Bvdsi4D
6U9sxeHIUEQsRvsmVp8ldyrUXNiSAt6Z9xisA+c6VCzmsshR5SEiZ2DycRHMKkfM+MN+4NprxHk8
Oe8JQnqTv/S9/IDAkdqPq6kwyPk06GoR7w7ei9zHBgW2brNm53kBTz3FAwDKBWBu8TJYnAmh3LV1
nfZ7meymZqjUueSkNGn0duw1mCSch9kb8FYsl5MJ7bFLTg1fIzeOikXYDE2Kx5lLZgVWLiOfe2hd
vFQYcDYpd/yy3FNnafdu+3ZceA/UK7gSgQfZdV+YJODC79xBAivBk379kigQzw/obOHRGjOYKkpP
v7TCSzs4EKQDJbGAhGr/yEB2Lg3UUVW5Gc7wLpdIEpqGRXJqW3s8YqFp74pnAErwVltBEeOIriqw
s7XmiS/izYAQUrDoBGfgP4nRQAwrChCzL18fjhHzCKCIKQTTLeZCTFUNkxnyPJMHyK1zFRq3Qn1p
TpiffBiCPydcxZaFJt/gXYKaT3eatiTMEv0UtZQ2a2D/USgKXZBRCKKZm6QuRza7g7fvNKMZC2xK
uTvXVpcHvypDfLJYImQKiERga3iLb1WffJ0UeAxOBSwZqA2QZORxErvOP9XzjA4vnqVYhONsyMrK
GINQUXVxSYOcRwr6GIKM0DnF+CBqD81QQ9PSjJljcin8Ed2t/JJ9f/yG9Lr8h5JTzgVThQB+gcIL
RVojSmhycAfg+H9If0yrBvuRgnQF+bbmyOorKk8qUL1KM5wO2jWyXoVJpDIW/ERuRIUepT3yJPn6
AmAxSmtAxH/sZC+srEds7M/Eyk9SQFtr4ggkdv9UIGQoDYwaa3B+GH3eksxz55zTOBRXXr3IPnVR
MOlFQMI3w9VxiCpruNNEzBHiyfhqADYWGFLZkmvq0uIujo8ylbNONAcOaY2FSkuBGgMyElasoGQF
NMqsqU5XE3AKU35aMAW2bkCAksQ80mwmE7XSUzf9uJ5BreDBvvKBeqvNZKLXxQP/d7NXuBaYQXpJ
+CPB3P823c0SpDydRgvseLnNcPSlvoaL3SJ2BkkD27IXuJ+nNBRG2lmsrkW0B1J9A352/KGHw56Y
mUTDiJa6VR75Q0V8ndxq/eXc0JTa6DVkHU1FshezqU6X7g7wmIARSkmoiNN5RJttkxpL2H1qsrxu
I/KSeX1C9I7Q3pIyxrw7suL7nKPOBGpJcvML05+dOI/iXxw2H1t+Bb80LLzNof9tufROrt5ffjI6
iYjwsj72c5l23BwODG4760y0EDsXOlv6aOeRYZAirGaQ0VrInnvcZxghLT7vUYBtfzPiEDvnA96s
nqOBUotBWVCouXZkm2qCNWJRaLwA2tCFAf37Qtuz4n056nD2GSxiqFm4c+O5oW1pcAeaVfC0fwyH
bJcFGN1qO8vNWgIcfBHNYmE/JgGq4E8oLx/k3J4kpsQ4PKDSXfh6GemoR5RFDgR6BkbpMMAMyM8e
tbvydbiMwupxjxexXuCV3sKi274K5eeCM30aeFonTCns8xNNoo4L4soJBKyCWe2zLuyh+/IN6bh+
9AKjvAa08X3WkCVsnz88i6uae6LWYPBEqtaE1oDARViD8jDzrUMbFm7a9LKwK2ZgN13k/kRY/6QH
ipkIJMCCA/ARessFcElms8Vw215dQvqXRKFsIN3Gh+M+rCz1RcmZBYFsANdFMaup/EvAwn4oH1Ay
TksG7muEryJQm+ftlBvwo9Hn8W/IOJb+mrjWsQnYHzi+sM87bZZ/t0gAUza8bbSvFVoX4163jgpW
RL4MEnaoiYpTenZooB0RAwWwBHD2zRWc1ObJg2PvEm8y1tUiVdoy6ypcJX2hcOnXUJnzJh/HGlf2
zg/lseLJZWoggOo6JCVGVblWcKV3Uf0N0S7BHDqH0zvGRVPuWlTmWXZTaS1ceMSU/0balAblnCE8
Clh3zZNvZPatD3RRkdRlz2lCmHo3VF/G1wbcW60hapGD8pJt/rG2cN8Qok2K9gai3AD01I7+60Tf
Y4oLcErivZc+nBTbwHvnY35m5eRlYWabbhoTokGX+3B0IoPfRU5TJMtC0qAZ+p3Yi90+5odZmcJT
//qNjfz1EsNHGKnG/gnJI7sxDWfL6WSV27BJtwqYhs/+31WrrWX21wXheYJroel3zJz10lHEzlxg
KUen0eqIOdlgBAq5nggkVS1lHxCMZYCX+ipGQlK8vhVlV0wMXYoMsOtSiZG/+JwIYaZITAV+cCEf
PzCNJNN3kKdNRCVnWOTa47bmqYauK2nG1CbbEQBfGIg4EixQ71YBuZQ4Bv5c78mA+WFlCNPxTiNr
8mut+4f695xd3IFNie46aIEXeXAmGUlwQwuKYIeihHlI2zMmEik8snQ4jPTqusq1lNFxX0oN3XKu
0K/KlAntcg2h8ECHr4z0hIVxoJ4DCE+hDNPdbUUcZfLE0ea55qcBoNy+R7TSeGGh6btIjzt2znja
agVX5+UuteGfCqqwP5JjvG3bFoROdXtnitO1iWlWxjh6f++bK6W6d2C11EBhHE+W+EZ5UJOfa9+6
us9YvHG5c39eJbWgPMRmkkbyPTSqmDyrg6Q7KGjxCYscdOkN2NHnptCmfRJys6QNMK21oJiQ05+o
W4EwX2Y2lnDosjHqNrYsBr5nf7Xspwk8WZd1Y+NkGDxMw18SXhedJsX7JbeqwIk++RP5Foaj/LE4
hoYPGCzhJfPBqaUeGlgCOYB2bsco1TMM91iH2cTu0UhJpUKEjRzepF7v9+uhja34oCueckp6bVxT
JHxvNRp5o7hJOmkWzYPH7rpYKGTor+bpiigHrUSQvo+iT0E6RZ9tX8IOId4V9ydIE/07IXI/Cpsz
70on3aJukCTiaLqAsIOkgfCPC63pWIuM2vBS8jLbVTN0WZq9/+8ou5XgUUQqIUoc1crexCe2fbuZ
wCQSr2v27SddJ5NwMsaGWb6bsIn6B+PiRBRNwe/yfN8oXre42dKgsociyg51f0c7Fwhr5EdFs2zo
KdpX7ONnIQ43sh9CUhAyRrtzxlcdREOftOiiDoQj3DcNL/aRNnHVcM0dvyhRjc2K9NZoRe+hlHDf
2uGrN0xS243FBziqF9bZ/N/ylgAk7sbB0UCKOvLuPuFDr6gniQ1bk889ysYVB49aexEh7dey9vuW
9jeRch4r5ZJ66Cit8uvOfWHh6KI6yfCq9/miFffRdpug+42BHmH8KuQbaa2VmH/4KtvwNlDc9P2/
qvbSYSKJ8bOvghCAojYHRgaeDf89npg7q/sXYo570q6ESYeirz9OhHQCYO+D0gdFsnKx8hJRtEgS
I9UtlNN6YjqKLuGVH8kotUDoIraTYckl+lehqGO9OfYHQY1QE08UjIoQPvXwzR3JJCNZ/2a1J+bE
mZCOkvZNYcwZwQv+DG01vmtnYkYMLl6C5C/EyAvhc3gL3bN7N5yuuqjnVUnUO2xSgB/2oO989Heo
Q47B7JljU4w7ZAnRIn6lxs5/8No+g5v1uff0XCPatKb0uQhj0dmrmXTzHSnvJ8zw0kFBDD/WanGZ
pb4xgNJ2rsjwt1wZ7AKcuHjeahkcz4ZCQsYgO4nqOn+7EuUJraxhgJMz9unI/AVDvC1O+LlLGvaP
42xPelTjdYVb/FBxS/It9l77q8BEk7fP7B80Qdt5jRM8wLA0ZDMzpGTOrOh7jOy3gs6LMvnYeA36
9hYepITYof29zGgUpILRIXpX9wvPkQtegwOsgVHyaDvVsK9y5zDATl6pVp+4H7Fh6Gi3FlUeVpG2
54SDD3Q9rlCv6eZPeqir7XWl4YukBaeYAggHvF6YsiwPJ/i/clZ/KV1w/xDixWjhq7+ISBMh8xOR
HHZbvcZaKrhbuFvj0/ZL52VX4ix1b4TnLD3GssfhiOzoUok/tkccjeEIwBo3CaFM1ebV1TGaLLAD
doKgnvISV+d1ya8EBMYq6LavJjY46A3BvzE2tGgis/aUJ7LHLgqXpR8Y1Puh7C7xPN6pbLxjjjMJ
omEZghn5lhaYtKF4Vs0fjgFsAwYZC7frxhxAToVK3jgHaivtK3zTbXFZg2+NdqRXnhS674V8ZiZT
I3j2MAad1bpqk8NEtAc/Gewd941b9pp4mg0dlVpdmPpwBP5Wmay77bnRhYi72KCVmSlulcBEQlv2
CBAtsv+nKW9Wb2dZ4NntvTeBxtVTpL1AaS2KY4ZBKFDXHxH7N1eknyqyssufamdJfyvFjzzbTVcC
RTI5cHKQW1lcfkeqxuvH8hXQqFFbyIbfqkFiq2Gdz2LANVA6kQnDjICaIDmgfqlcdBqFvhfB0zgG
7ZGm4a/yv12CamH095jDKawfxnMD+ekLQy01hAy6vej9oAEvu3+30CSy6gZ76lW1A5Y+YYnd/las
n43xXhpWhEL5M63PipXxSfkLIHt0jWZgk59CD9frP4vTtUvTEAwQ6eK4edXvvefRzjMlv4n4f1kO
EH/j4JOSVCDZR8WjewhRgp6d6otPYT+kvVaK4hIeClxY9Nx7Cw4LtqrdFCIzF6h2GzFxinK7wlvR
GABEH0FtAmIRpYrZdF3AasvukGt/UhxRbf1J76KI61M5oaLr3a3L7FlTRoHbaiNqZh07yAce5seS
tZ11SKfCI/Ile/OQVQ3OqidyDcp47FJxMKmcjvIS8N8AD85U384BpGM3hLGTpMzzkG+Khx3UEQCi
l9xueiPd1ZmF7pt0p199Rc44KCmSfBj9zs4Nw9p/elCnjH/SFnnvV9arOUrFDZsxbB8VMgX9ez2J
jeHwuYmUPGM61IMi3+fCiMHbCILZbMdTf8t5/hjnOghXHt1IBTVpFkeiSUkgKl5ZpxMH4r5wz8To
I3HNIjH5E53Z7W5gVpvG4bdg5QrlgHkI1x958b+XW9XRNRPFiXfuYzKF78YxrP+oOXc+trJqCyU0
mt3yi/mwjpMV4OZ5Bk0kmnDBXpROiLo9U7hL6uz/SEbSnXMPmNRkPRDlG7q1/YDQ5vVjXXBW4Lxx
vmNW36IejavWjdHsCYDFwPOVqZ3ew8eOubQFcW57478enxIT/i/2lZPp3Yh/axrLYXP6Ly8fqijL
Y2+ejD5kJxUB7OScled7NYblaxmo4xk0VXj69HIvF2djkVV+uWpWM2Iin0A0tZN0Kds8AL0rh2gn
cXs4RbJC+Uxt4tRIo46I+qCPo79SBjEdWhY7Y+I27lkjCxywiEAC1qZ/MaxzpcPJCejhykZ0oDmf
MrWlndNyHAGjBIy3whQ8ZExUCNKqUCU9ZgQwOGxROkFXMTchv5T9ezycoRdy2DS441b5ZNJMQ373
RT6P3sYcIfUotlijnVIrQcqdiIkG/H/cZ/fbiReso2w/SxnFCWkbnZR+c4XBPqAjo6e5Nhe8eDyO
FNOzVSUoc+G5C4GZ627soTylOuh0AXscSiyDrQXAvwFQ2a3JoqJ6sJMLT1IM59+oUgOSfVRMpFHJ
ZtLrtQrMpycrHWkA5MgqItFtq35i5YTuuPymfWfxRZex/ZDdS/J4v9WpqKqx6/gZC+z7n21k1vuO
sS/syWvn7+u5bltCVrii9XxzPGumpZOmxOCcDgpjamhndnIZYRNRLQsbdR8QWQlulqh4J6O5rVxI
lzbAMl5yiyz5Gt3rS5il+n8EbsGgoKn7drm1zhOrgngOlkYYdyFlWd0BAyYf8nnS6NSQF44gKIb5
8SAjABTiR8ysSd1zt7i87JfS1oHOBpwHLcl0JIk4+EaVyc+Tmm0WwCbYvg3z3niR/G7524PAdUhj
Kcp9XqYW3O+aQX+WSvzp/8fPOoLz5m+yYDBlshvLDEsuEayVRjAW69Y92ncifVKtpWJJn1c7eOd6
5vr7FdMbPTqGK/5oSaM5xLvrKp5Vnm8LHQmRniUvDD7B5Web3xV0OnoO7X71EYDt6aTeCgb+aVwe
65IDN9Zj6bsWJjh4Gn2+S6niK+rUbJABlGPDa8ycvwuhj3udHYCnYrzGiFdlM178tyBSVCKa1Tj6
K6tIm04oFFjq9WB3RpHDHO7Hc6Ou1AQ2URI39dN6tTDp5dQPljXVpDUfp6K7eY/40kpCS+U1ufpX
Zg0y+cTvlS4oU0GJt5/JJD9HLKBahF7TsL6/QcXDXGevJzF/nVUboZDqUeE8Vw6KezqsqJb622sW
svP8+sJvs5SR6cBvtsR2LW/T8iGOrt23n3JoAvCbCq7ao91gBm8ucbgSB84vjVrLK2n6PPdL9MoV
ZQubH+bjBZM6Ox0ab1Nauz+uvXMZfWLRsVSatrdUuvQNr94hXqAi4DwOGS5U0Re78T6mHAMMMrGc
gOO85jNLyuy6oXrKQK2izMHM1785+PNwDeEXnQRkO6AqcuhvchC/+hXozq5kPyJqBLZJCshmeyOZ
5PWVCAaoVklBivGdkdO8sIugzYHBX3tmCcpO2Dklomqfy0utoHZRVZi6mHjCUXK3/x2i/t10ldiE
+sACZM36z+EOwih3y9Fz/j9ynYkgfmvsv8+VS2KfUyEsANLOAa8KNTEfE9OF3h70gUpqe0La9BZX
dn4Wh52vyzab/7tFj4WDvlY7MEmOI98UUkSLhC839yPREUnEJd7CnlChsQLbqtadKQgSNKykMzf/
IydEMBGVzSP+AwxlmMkBH360LPMVpoInulMyZ1MkAy+E6EcUYOsKieC6i6MLvkQRQMHl2gQsiVbo
JA+XPQc3tcntFbkOfBa5clgt+QRmyKAy9pKXMhDjs3gRzrv4hryJJoUKPJ0ahSUX+tyWqWJzPFmv
vZ2H+OZ1E16u8AlYuuU/OC4K1Mefc8ZsgtC3NC5x3+THMiAysdS8ZJgDrNnn/mUmU7UDWawPXlxI
t5rgWQ6BM77u0n93inL5imrMWQkXsDoWioDpFAUI0rlj4vlti0EAs8UiHXri09SNoepzYP9/wDSq
zAVE+a3dsDcSbAmnph4JuVLwi3E1VDXNszCcmQYI697QJeeIOt3x6Cu5pGrSJSmDvCwvqlv+XEHz
lyZNoASwioTe+sK5C/bRPPQNSio0HrplVx+Jeq81DniDIa7MYrpcJcCOGpujcKKp4c1QNllwNKY2
m3Sfzh9+P+8NoSDBGGvzRgvbloUa5Me61CPCSJQcTT90hkqT0AmoCi7FDZzc2e4dQK/eh+St8pjn
JlljKsvbmL/+VgF2FeqkC6VWNxG6RUZuzpj9pbhOkqQHg3zKCLObVQ0LuhA9LemJhEN7qBoc0zvr
0CTVoZxMtM95FnW2xHESMgefbF7Yn46h1htFNvwd2tRW8yYouKLDXJp0WTFh5w9aplTv1+kEUQcb
6MGBzKAM7krZ3PoOY+qOfsWMXOPbf2Xn5loEROTOoPXjtbJzMUL7QQ7uWcT0H9jYWyOpoNVByRRc
EhDBGz8CdKc/pOtCXr8MixuuL5Uw7AEfgcLhcor0YkDrYZUrsWZcu1chskcuDia03lINub9P1OYM
TuXNyHxdHRtYlMSolSJcnNmuJseUdhCZ6LKt/pkWmvMJY0vkRQ0f7LTCyZuxSpAFfaWB2rMiqOW+
0fHh17QCP2+aGw23p06OFYKhTlvkdDtLN8GnX90inOKr5OqbhYC0Ip0Tzpkq15tEJk1eQHNXnkPV
SvJ9GU5HGCeS9Hi30YrZOkLNV8FtIdOyeqz+bfrzhBt5G9fK89CBJudtxYC6M0LFEzabU81kGIzZ
46sCYBFBhFY0SyC8MaFY8x2tvfwKzfXhACQP9EPtg0sTOC4NRuA/8WxHRoxQySegPETGT5sztaFK
I8LqY5SQXfPJDGwfkU6nYfJaXcg0nzYK1o3cryWkuyj/OrBre2h6S4pQhq8G40+ZrjQpYzUfVNAI
hA7fDw3kDPO/xgNW6rVpaiJM43LHejpGfiKGF0716zjNeGHdXvW2rwD4fBdCHzc5M06BYyWqCXva
n32/qYcstnypXuRi9AGc/Wgu4fHH+/s2d80mZxysW0rnxKbUpcQ4M7Quo1MA8yGHy8W5Uebb4Tid
e9BD7v3YVp5U7fNDH5GLFafGTDudfqcAOfEVdM/c9yFoGvMHGLI/yQ+nQZrQfeMqQk1pqlSBOj9P
q69fsmeIFnxM3vZK22nnnC8UYL0WaR+0WDmSJI/YgR0rEpVNwcOZ+M9miU1f5jxxi9Ydn7WOlfD0
xr3osoGyZUsccUguEyCzUZCeJJ9g0EN00nB/xO5LeCfv9Ni+1NlaNXibJhuoZrh2EZL7rRC0u4aW
2uQmvSvjfxn8axrPasoMQDQ6FLc11UTjjwssw1dU+9lRB8kWIwSxdkNLZGg0WNQYJ7CeNeuPIWwk
a6znoUwW9SZoT3nvjer1/ArDY/gpt5TpGP2Xlm+msxIIP1ITGbWIjwaX1E0pcix18v5pfPpGYMSH
OymNWTxKhnbU+Jh5yDWHsIG/GW+f93kVwqomRiWDChDW+fsDz8KvJKE5wpZ4JIPQjnjIkuMKVQ28
rkOpTFw3YvnF0OP/+V0yqIAYKHiZYTP4ow6IVf7rg0z8HsJFCxNIwtB1FkoPQlI1e1GZZVQT2KFN
6HqwgP0TYK3KJ3QPupQcXCYWX46Peoe/FIAH8TFWlGZPSlZAOATKZj/xqct31yHNUqWObzAXOcI1
hH3iMlqJ3ZhK+G2MXGRB07ATxyAfgNEGeAyhtXMJJOm1EmkApVuFb1D3enZoqpyYs3nhkkXsdbSb
vmyhR/QLr7mULcA4fLfMK2ThvXNvSodyizabXlE3slzZlErDvTAfjQ8c+VKtz9q+L1KwX5EZ0DVP
Yes6vU7iqEbjjNWFNuM/pRBpiYBmkfIGF/y0Su6soImxv9DhfU4m/dVSFejjkhWd8qyY7gEEVnc3
FGlclR6Eg3rXj9keGcx/4sgUzhK32WI2bGM0pEJWqUrfJeb1pygJr6i8L8Cq4RaMRAlMfam+oSLl
Pf+uJJbElGmqSAFN+Q37IOlj9oDM6STKo8j+Y2A1Whe78ZVjpCzeCuIMqPyB8KbB9cg3vZzQBoXl
S7LAT0NyJaFApWOu3FHQzbCgFzg272SrtK4W2RoCQULOG3zHiJmZs5l88aU7Hv+DE+GwTUvofFkq
0q3w7PRngh4I6TIrvW31SlW1eEz6SFLld4MZFeMZAu7+ktSnQQL2tD+EDFjbW5oZsvb9yAnOLsUH
24mAawr9f3H8nZz2XXkwMrbTLXGWpKGDVGHxFnRpDXJZp4JxNDZFbUicYxR540OVa18K4rXeXr0U
gsMMprbEwfWvEJbDzajOEjgP/SxZ38z1/ML62aiD3Dq4QWw1UWnHXf0oE811td46mxh/8SJ1QvyO
DgtN2P7jkAFqJ7g3Zcbcxws+mynAvIi/p8uQWqGCJF+w3kMtET+PxZ48HOWbJCPLxERTfdfcVYvJ
MMaeBhuLXOWrdjthAXCnsFNhPP9t8vdtreoqmz4UGeTNs7HQFL9bTjQSx9hzyOkJJRA5UCBIo3l5
kAqYY+ZaI3as0SVlgozcy8haBO+uHGX4hFJ4dEWVbj3Gj4rQK+BsmEOwM4PSCr25Utt73Whk7Js8
ydMZPk6WMY4Vn/EriCioOXKypRlkzuT0A9aFVPyskjYzUGCJK+dIc7itHQFLER5P2YiKfq908RZt
U9BdMqITl4o5Q4gMShtdTsIlUZlhyb/emolo1ZplBAtU7YMiRyrdC0Nbn+ZpZaqKCr3g/tz0Mt1i
uWbHjIIwu58du7MRt+vCqZ7crJlocGIUamQpgxV06WKR45YI5ImJJQD2odal762wm/IdW5Kl1hOX
SGfwCLQUqVwUPCHAAgCnwqqxlQd999HEJ3qF0wdcO75cldhaJhKK2wLMWRq+8pd6t+r+F8N67QoV
p532qOFMPocbTGp63JckDC4+/eW3B+YODIyaBzo6WuXD2vUJiS7PyaUdkmGX7SK37OIhhxy+7UN7
dsH+E2pcuSQ4dZM0XXWqYoFd6tAsVs2A1BAntiWLUceqV8zGA2UDlwRzeODcb2uyUlxHbp9ZloNn
iZgvk0rxRMaQLpRLpCA1yrEXmd9vXs+oit0f8Cbv6fRYEaUF0Xh764bzLIzHnb7oqmvv0yyFy1g5
4gfa/LXHPp7GezCQMczsaGHhvGs9HozUeh+Gc726S6exceWEPc8e5EeIqfUDdHeqROLqF5ibkh7A
TjdsUVMf35L7WisXaacMC+8DXWV+UPI+68bB1+heek5vadh4F1A50fPCyhScMY61VRFhVyAnxNAC
v/Y0Sui8kCkPueREs9HAcPxqRoZncd7MHnp8z77+od3YZXMcOYeH98dUa4N6tQ4+HZNawoG62GCk
JTEk5CQv/kbaURis6Z3wM4eYELBzGZ+g1VRGnfff52SQXSC3BWDL05oQ0+6ffpi0AmNCg6i67NJm
An9LXXURuLdLu06Gyk9ek/9aY14TlzKBdE5NInp/X4YMAJALbwqVHQeenL8U1TM19Pe5qu399/oF
11njNWS6VhVnIBoTXKQ0Vg+1b1nCgUeA6fFv3CIyzAy9dArN03DRP+P2YgSoRjfQJrZaCh1iep2+
BSe0u1aPZyRETFeoWQxTvM9sABGAFrrallDMD6Q8iJKjNJAtPrqUkerJAF9Sv4U11nj8KY5/Lj4a
nnZ/gFLjQg9mPB/+MWZ68bvPcTfjcEZmfoS+g1qAlmmkUb//f5bg8NMztKMOfNovxs6acCit8Fpw
s3LehpfGoZIXARiAVE0HbznxAK2WtfARxSVHZPruf88zNbB0jknqZmejJGsSVrKgEX4E38xKSFKA
yF2HH6kIGIGEP0fgTisAvyKyLuusJZT4BKu1MnFkM46Jf8eR8/YjOp0gkxk6w3Gx2SV3P3NY6CfG
6lnxLwXVd4ixQejt4VppZECXMxr4PPLE0utEoJzj0MCWn57+3HQZx+p5tZ2KlnwK23wehf7IgZ+M
3I8/Zz9CsY+VIW+TulxmIhzgEhVBng47U4WN78EDT9GfRIVXAUcqZt7IaOx9hUQd+j43NL8O0moX
PuCyv3Z8COiDY3xy7YoLAW6dOa4fLz0S+fqbR9SaUUHHsNABfzgmZHgKxSwFOtY2OssZTObfS8MS
39NeAOOKfROaXO2yKPFh55osjC195H/jX5HbOOfAg53HLQ8kXRq2nWgaEoab+2laFMvD95gylKJf
FworrithjbJ+p0RxqtcbFUT7mtt4ltd671HQ73lnuRaD8AhFVCKEj6Gu8YaYBz3CnZ9nxPdnMqWM
Q9l/2YK8fWraytVZ4nNZIRiTrQb/1boVF/9/r4R0YlZxTG16RenaHPcCHIsi689yLG7204yq0q6U
OQEWlLHfvoa31RtZHSGqOi/PUO99sWF8qe2fcuCegXBjuxQ09IBp/PhdHrCRA1UypTxLhgbVwc0e
XFrLoJUi+KNvO3sJDMyESm3VBo7seVyC2dxstyrdb1nYckusdanVUXy6jNnsBbb1ewpfIwXLHT/A
lnUXcjCpU/JgbVX9bPNPSvjvpIt37fxdUCdQb0nierALz0uPGmiUuhn5C3oWhsKPEl9NFbOQK4UW
GcjZh2U5jEjMUb9G00/ptfIVr7CITUKwZsWTMNDneawWp12BaT5q+V+tEDoO15D9Gm1EBe/Y8yFq
UP9DdJaG4ce2+fyr8T34lTaVvPUPnILUSAbfCWBUq79setOkVWtm8vVxfdmgahcSvwfSC6VqjheC
DtvECk3dND9UO/QNXzdN3Tk3MhGiwH80TfRD2yCT6NF8vD6LwXQXgOAiknUlVWbV3IRQqivgML8F
ViwRrxIwHLpZV9pnvspojYGrIUnaGUarCcWVme+XVZWlLkOiKe+WOqYfXCE0+dI4OQ9WGsB3BIBh
gO/yetqdFQHLAEw96Ld/L9BnW+IGxNqpAyMei7ebocZ4e5PaKWwsZcbEBjzcSDT86hYWK4RpEq0Y
VVHc28NKPp02iuFlUti6+VuvuNa+FYNX2XtqkNSY8Yur4Z/R3T/PLKnGib4zgn/r8ekDZTz+bFGL
9ZCFpcw1gsVrgKmWdBYEMYhXVFm7H44CC9OqxmqH5NEdR3oJoIrZpx5ml2jkWnei2idDvHex9wCF
Bh6R55NN0d3SdfaFf5UPj8YK9DJvbHG1iM0YvaQJqavWoYX2CxXSGZls9xAW9ho8VRCt/HqYp0eB
lMUr/eG+Yd7JOpmN0797NvRoYikM+/cQhOuCI2kkW03cUeHvTu+E3hwIbamjLv/kGj95WFsB25rr
xoZVk8M2AtillHK38wIFDwe40hF3JIPKbcyWEE8PkUZ5MCWDCHfPApQTvjT7DWHoO+XCG6Wwb5Ek
ilBufIToPQuOR/IqSDAINnFQPFUjXrUCygpTeyNDZ4JyUF0N9/a+ccnSIbhnVs7tiWWJ2zIWg2Pq
+Vf5y4BZHsp/c+/Y5PcatOL4p6jL9HlxOTnLAxaeQkS4Yh+tC+/xh/jarA2EI4pLalcvZn5QyD1l
eywkVPOyAhNzaL0G+luw2ct9EXu7cgE5FrDfW8Q4+t9YJ8uRdKxwrZam4D0Nbg5ZQ9mqNOg/s0xr
MR4E2ehfFWs8gfAZYzdcgi1Nsz4EZtTYtDqA86O48jmmJ2efqvEoXof3UDf80QXlEND0uFyGVgpO
2hkTQ4f5fSI2dIrigJLKBGRvzyxQd2BxbrykIkv+JetgnJo+dR7WAFiMYDtQUJ5XlHk7T8O4qWn3
5WnL5j/SHIxfkkRhF52b88BYKPVAjEx7Vf8YuGuQHue/e6SN+qtg0PXCImyZnoDzQyNK8a3PV93L
0QFoGVALPPlYKLG0H+nCS3UrZ8BWh/bSa2h5oB5vypchxnGDjzGHzXqCRIdcXjRkFKuMcWuUKhVV
LoE6/LFN349FQ4SzNGxZHE4nhkwj5RRKcrb+JoxUPklqi2m6y7IC5aPQgoep3t8Lbi1eQ/ZrOgKb
88R07TRdjdDcEEJ70hXY/3jwrVRQpj+qaJhsNUDwu2aDtiMl+Lp+ElzT5IYHyP0nVfAHNaxu5ZaA
LoFhrZit1d4g5YV9CgVU0SzzNo1GCUmSXZBdEsaKsGcH6kxZFNC4ULKuFXdLNFnTuf+IBXgQPlLt
kShcuufSP1mZK+N8GC555uxvF1N0owF/8CKfhCzIK3WolEqWe8gqDLKH4/hJaz4G7TzQqZ4r5XQS
czdZObloj7EQXa2UHhXoShLEPIg3tI6JQS5Mkb7ULUVPuW8peh4HTsIAZstvFKNQ0zqdS9EWMx6J
jBAynZP4RsDwmL3JhDHjml5a81a0ry2WYakUcMoe4wVigYVjI4P0XeB+k9A+Za1xWIjauwlSzI6U
YDLcD5zEpwKw5YpDsZu317TwMQFwLYzESX/xK3bVKyXt3I9qEm8OM93kEQHTSZ+NYPT0y6gvuSPW
44qvmNKuGErYxg2BNYdbPhx0ZhuQ/E+zz4zdckKoNupCCF8pASFic0NHGQSRk9ogQb6MftXb34kT
D1PBcB+GoZmDj0A2bzDle2QFkYTxrPPlh1ueleboPibhZ9SBjrQL+rdK4cV6TqG/WrIBf1yd9Siy
u4wb7Y2Tbvj1XbIB8FShe6RQBv4ND/M+I7wKJZjSJfWd3x0OfrV0xPf40KDeN5jRBn+YrQ4PDraN
YN4+Re71eyshVuopeKj7kqhppMrMSavtgRiGA0YbIqhH5XnBLKzoPDa7lz+bO/C7SUPtZfSHtfA7
D+9aYuZp2AvlNAPKK4fRFBNbw5/rR134mVg1x8Ho8nZDZIhQsG/XGKKaQ58oI9ZUVBaVAT0p11Xl
cZBwgRLwlaneu+yfZNVMUwEyfD/8xMj9ZCHv/7NqTK25KWGqixS4gfQgGjJeZE9RuVQmgiaTLqHc
pUWi9VsLMR4+ao4PJKDT2GDa63VnVkFuSDFbvy+/OKZg6Sp+Evhc0CBqM1hjpFb9Ox8Vj0bdrjhf
wgs6/hxzISIYZIZFDM6oj3fhKOYE8Kf8+h8rg6ZYzu3hK+h1gRTL6+jBJogDs1gLH89DzRVT1QiE
+Ec2rd6T85+X8mTYv26ZAp4ndRMrFiIDwoEXMd2sBg3x5+lCxU+yNl0udm7MgGBBzuZTR+iAcUNd
72EKjL5lCRGT96Zl+ZYKw1lstiaS74Qr5aC84ue5J9JAoHjFI+pJglmBaxuxM70MRwy0cdLKJnh1
F92umTbpnqvakN2OFvqiP0FU7cWiPW1eiRoWdWUf5495VHHjKudFFmlJs9vpDKmrT5Q3UhERunWG
NGvLfWRBc/+3S00m7X9jFYudGnqSt3k5WcxiUaDhT1gaolEeAoG4p5nW7QWDk5UW/ShkZIqEoFG5
N1bV44U7xtAFww88O0t2blPXbFC32sc7aRqk5DoBATZEpr9eu7Ot8tSNKTqKDljYuVZwBVIYv1qc
ZITT3MFAD1VmKBi0mKZeOU8r/lTGiv/GmNda5Z5lRh43QuUfFvTEqetjgVCEgm446jCYhW8R5x5m
own4Auel2Qht/jxDnqAox10OMfCgFiCh+821+UXpIlS0XzV+zB/lLTxpPTeBj9ES9fgsjAsHwi1c
fdDaPHLfgLq+NE/0BsRxYwfzfu6M00UARaM8BvuJc4yEx57JrppXUau7KJQWHFDpzcCL2ILrT+R5
tuRkEy2qXV3OmbN6+ue/TbW5nd0CvEuIvyZTjgf7GVd0ZdOl7EuMN6vwF45qPXc11dJwYzmt6PDa
PQ1ZPwO67zozhx3upzH5ZsWV4QHNqasF5DjSWBQ3YCJeD1D4PoTmGvEKt2GevEWXkJxwFUnd1/hz
BBwFqExvEI2wEH/4zkyiWfCid7Qzzgu7np0C7wLkLFJuDAw/FhvkkOWvIGn3X+8tPO2pB5yKilA7
HJ2SrAXNemStzHMXTHBZ0bNV79PfvwK68HSv+nLSBX3ynHzpOd03pCA+n14nz6m4Cq+/uU428kEB
GizLuuLz7DmTjO3Vvmi+uR49tv2q5cBbQlXaIg7bUtb1jQnlX0dGUCruVcLeg2cP2yenH3H8EaPU
peOCaXvrmLLpPLdU1GpEaFhCjpX3bpDQdfn7YDjcYaWIf4PHzOolc+uMf/UAcQGRVfJ6p7SrGkGu
v46wfU4Kxo+a5jzdKR5LF7ROs3v+EViV8IdxMnXOIb9E8wbPw7SIO41ghEydhGGrgRPuQc9lVd+2
iok0i2mbdCYt9/GVqKOJEIOIR8HceDoJ9EMNOgJQgQ+eBxjtew1ccngE3Qcyzccw9zyt0aDS5rVm
XOf5xADNNOb5s+85lC0ciIkz5Z0sFKd+sEcV5/18ro8RIfVU8T68T4J3HYy4uzswtnLRhtCih3+T
X06E06Yg2++SYvvS3hGeD11EEr1X6Hf2T/GlF0PVwV7vCWJ6SjL5suHebEaPeulrx2aSzG8zygmG
NyQZPUCSQuVAu25b0K0StBENB1PpVE0X4dH0S7xoJYEI5LVglAGJ6P9L0yPO2OzNXIrExcVV2x9a
H1HqnkMz3sAJl40yv30z66bh+MgpSp+rUZ8dUwjeIpNX9rNoQZK14+ci0jUhFXIX728fOw5e5Plb
2oIe5rX3uRhhA10vh7PdwoUzHuI+4/d0whPSBxrMLHb1Q+U3ZMWG7Ft7o1EtAIwpMXR/rmqCqyZ5
AJ7DJbqHFonoTLetjO7KQ3SIN4HBzLp47/QUdu9SjyEyLSQvy1/F2w30wOv/BkH4WvAfRH71uxac
NB33tKc1eiK40C/QtuBw92PqNOL6rb3KC+Gg3yIgqdotlKqkOYrjlFxsBNJslnjG677ThHFluuky
+SQWtK1Ld+4MPJ+Bq5p2cIjab8GsBGLKfMXVPVtUYFGjJwk7TcPdgmWBoJY5PqErl1/WUlbjc75U
uytmlxEO+WGnZLoHb9f5XFqvbIP8eRsVl6ZSBIuIVYwUy8bW7HjooTE+xT3Ruq9qWCkJpxjOq5Ca
Xqz7ONpzq+79iFiDCLnaAvqC6y5oSFESOYZfyXabcZqe/+DaU4wUvrHLkirwFLRwxQrNLAd5h8NV
vMRsZbu8OFXTv3dRRpUXZfXlzgQP9ua9iqEqWI62NEdUspXLK6FscIlVFPS0SNZDSPevWjb3+6a/
R3vu/7mC5JakVRM9zoIW9R6MEJup3BfabEquk6g/rY9sSuPzK9Sv+y3iwvdW7PIMNv1ww5TSJkh6
Em+gvQyAqDVIoyRm7PlWBjLQ6UwJbWDiXrDcZxEw4j1gjZ+RJpJK0rD7z49acFQXaU/Ntq5eIJ6H
dwFFVr7MuANJpH8SEKkZkDlXqszjI/9x0arY9XG5pfRT1OP28YRr7iCT2FJw0BKnBEJdcve4bnsd
d/80GZKlFxuseID2nvCHYnGVirn5i9cPvMJEskBojof5qyxo7VRbWqW6wuhd5Hj35K4RxOgsi/kt
HK2OaTGYhnPbd+fc/1YUMq/q0Fy1LDoFkF+aOFi3fe33hXpdDCVUYEs6kXc/NfgdBulARdDhOgsh
geENmOL0RorlBDDEDsxJoTrgFzYkE/SFFAwnlNWVmZybvk5BB9A5j+NUZSENC0NJRDPQ2oit4INO
XHkFC4c1Hae9GdABohXv34TTo96S93oImh34QKcZ6CxCknNKv21gNhJ3iYGPcOA0/JPzwpfvvbsT
YE6qBmtEi/bFWQ5nMJMhgGx29xFaLuNbW5GONxTRJt+3+PYCPdL6PLMzM1KPLLlxV4nOgm/+JuXA
hnUvcOd0VyL27SE/GdziocbAgQgBBlmusra+Q7qDzwLUWTQZvjt9pgekYTZAbZLVYhb/VgrgUgC0
qEAqQJrI89oQkX11OMebAuRXuYh8MfIHBtYuu3IOEY/5e4qP8Te575knpG+viPb2B5S6aCsx3KN3
HqSRO/ydAT7mNa70CnVefUbnWN6ofkOGhLQUE55/MqnjDkYi9iR5SL5LQu29PG6TNmPLN92fGqU+
8zSYn6U8p1+ZEW4jeP1KsdjifwJXzEjNiqRUZzGcJBtTsQWLSHoKxjxDg7fqHctPo9cJ4eaVy4oG
Qn8S6xqJtdyLmw8uei5c6dEVdxrix5/mMHdLbh9lRPPtFipzVrxkrflpZxSopP2GVZMr/GymCqQL
Fnvb6DpeEZWMfK/P69SD1aZgvNLfptaNMg2aqcj0ONsH0hAyDQDX6GDoBdRu6E6qiW6+AyiYWGfA
odEwKj5USzbL8R248Rz+aTJDedjQ/9wAqNqCPFkn3rO9fD8bwbH/NFzhXC3soAwHlQyKNX8Yy0+a
gmcXY6Pg3MnXce6oReZ2/HlUesW/lo74evmaXhVXVX5bIjKn859wbHmRWYdymK+6KlvHJLDCHxMh
OEvmAnlUjG4Zt5YYmAlt5Nq6awlbK2HaKX6+mBqx8/9/0lLV9nYHb0IHyf69mFNTIOAMmlNFodBo
tZO6+BErj3UAKUCQ5gs0dZ7G8lHuzHj5xGb7F23xdGI+w5wXMRlI3+Uj1/QtXwZZDQeDgh9PyvyT
MPuM6GaXFyL+Xja5gEaaeJS+F1R5tgE/HHFiOYgFL+dAlpJVJKpwHIxbw2nmnmxYzjGrY7H6C63A
dow8fs4EJZLcZKR2zZWP3QJ7dpun+xpEML4rSZmLK17AavQDebg4lKQ6py752FPExWse7j8OcfRn
/A/9kHDYMVRhXsr0bA5Xzo+9Gi6y2JS1RlZQRD8YPXVb22jy6euKv0i7pFuWQTl+QDUEbRELHMPD
gMcJJ83LEKrpcck4bE/HUfWVnB+283C2jiocUfaV5TQJasS0vlpHZliK0riG78SfpUSKpw9GsoxD
h9yPjHwNrJAJ5UiRvEsNGn4lG6UCgLPhUBryDoMGlK375nSRacVTx3HvI9soiCIKWWw1YH6P+iT0
MuH3MUWRGiddfJwgIijVSfPh2IMln8U6kHdFD5B7geyvasawa3Ct/mU8xhnfEMwAU7y/jwDr2kUc
qfJQokDP0aZO6/A9NxEFG8jh6xUaOf3/DOiNYl52hMUaKvz59gR/MnoicGM4IxOU/xl8HKkhaUlr
/lT7OAm04Qypj22Zycg1W9y9vMkhRz0i0JaNeXcRMJS1gDjAPWyPBEGnE1l0D07qGrRnIY1sejxt
YrWdPvlhezKcyanX55y7tnJa/1a+g+mRI1fye6WSYIA1qr1OXo7j8926qXPK5u+HCJLhMFKoz/Ii
Tn7mWXt4uYjym8jfSOdy3OMv4a7ZrqIuTu/ZwxmvRmaFV7YyS0ToD9WnzSoOlcxEdGHKnMAIV7fD
efCV98uRZlfO09O3nlEq+drpBSCqpDt/UvNGtuNCJ1P1mRNpHFk+4pIxdC7ZMHhMCo5goMyZQhUF
7bOq/ZinjwF0nFOPXvH6cYEpM9bJsn6kL4cUZZg/brcUitQ6MkDgRzqMUxR1mNT8FgtU53RD0ht5
spOt0UDTfU6+UCxQbE7Tts0QFZ/M5JRZauyftKxXlXmHi/8QByJ8oVhvgju37M4FdafQiRNYtUeM
YhfHahAz/dCFN4G6aQHHrq3yIi6s1GFxnxxagHPBIpPvgfrg+nCvo5Po1tZC+UOdjiAeOhTQiTxc
BxfTRckq2pda83eF+RBfMM4F8FrfatKkoulZhLt8zLpyTVbKzmH5FDu6O8+GM/Egx2yuAAqDiIg6
KPG1yKR7iUzeA/teaukw3dIQd7S4sOSloM962A0OilXNwUgjJSk4+Y2BaLX5XJEXO8fFp/11WsnA
S4aDMlXMY24AB+3OgT3/VKO20NqhnMeYcP+0ztYAWfdB1hNi17Oh+0DFBOngRtxd78YKuSH7sMBA
GlpF4ADG5x6r2meyo6kI5HT/Sa7I1deD3AFBkOvDkCGTc+h2ovnlgPNfy5EjmcR7Gfk4l9atNt4u
jiLksqAwBdICixBQ+uknvwUxqef62Ha85tMdPe2VUbmCKjZYb8nXSJ09GVX6XkK7nxTAY161FcLj
AV/G0v+R2ibL490kRXehm1wzxRr5Or7+GVe+/8CvBGRcIh2zo2/Ft9487yGaDnThEEyR8D0SBMQT
1XJYExu5HsVJ6yhVfMFxYClyrmOuHl6NzaQBSgR4e/e8bNqM8lPmUF1td5omo5i7T5jr/BAsLMO9
gnmDo2Ao8rLYyTuD6+OLyuqrj1W/NVaGkp1tbWyiplO9fzsNxZSFbNo3sCthBDY6Wak+qQKFidxg
XXJZM3uo/aboFMJvPMvmazqn6DdEH+6km+6RB5pj1Ghraqgxp9QryYyHgBYmKXeYzkLdj6j6YXIV
yrjRCn0mHeGkRHlHoKnyeIQtPu8ihyn6sQGRNJmxjOUl7kK3ddbrlHApl+bjD8anpLdeEXkTz2Nq
h4RE0fCsaUvkGKkraqN7sgTPAlDu3/cfM+CZGOk3z212l1ZadzTmEYfm1mb0BBPfJcVfM8hS3uAW
xWQZwbKM3ehqqGEPxuGPT04iRJprtEAkCHMgEE2sFSC6Rm3mSoIfsb/v9tMpHmBnG60TuJLFUBmf
Kp4Hl2CBixV9pfI0aXpwg/IeLM2irfTZiPEtKNP4vGQh+MgvCJfDaQBOFeM8cnXIu4v8QnZ9zWLy
M6I3v5S6zgDCkZm8JrwdRI/I0O8lWHgo3ucxI0fYjMSvc2TaLp4IAjsQjB8PIMMhjcEegDlDCW8r
yrpgMj512d0l29JG5S4WcELXvbLxaeMXBqFYkkT5ENRrijn7/+7lUGBeWhIkIA6R5kp8Dmw/rn9S
w5ZNxzpAvHlAFDrZzlg91hZ1oMpDKqivKU9l29UrWVa/si5GvblP49/sN2ND5lvDGniT+/U0ysF1
ZrboQtrKuCmKZQjUtL4PZm8o/CilpB7Awn3M4IVJ8qJY9NETWSrzmSSKa1I8El+uS0P1H20nelku
pxCU+lFEWun5Ko+bTl/wOh1RwPPtJOAHrgc7vvYkErJCvUs4ViOURqKb1i0b3Fr1pYqw+HumskBX
qlqHqTb60v0xhUzSP/F9fV+W8kJHvVatbnv+lH6DADDHDwPYU0pIjJteV591J25hN8peUzVrOOM3
UhEYIaXFB4dU1PZGhsyFFd0jcdNbDY5mdPCGa14ecpbROQMCm0+ZL7ygH3GCTkAsOeWlFPRab+gD
jJ6KSiF/vOqCbQ2LenkaMKATnrTC13gUjvqTjlFrcYPJ8byCP6/6PZVvu41t49ZhU5N6VA/ioMTI
6Fp/h+4KyV0hmJ4aULEFnOphjxRtytR6tyHytTveir/8tbhBbZzxv5/XmJ5tRrRfbdYVmoej5EdG
3Zb1pglEMW1DGO8MCSx7D1HvWgDgu91J8Z5pklc0ury017KjGWERY1n4Oc9D3R39+DPnwxNO0Y9N
zLHAuq2TseYTFlmmCPnwqJN7XgEeqxrg03dCKoOUQYEm6tVbu+K64N+K/KQk6WB+fuLaphUn3bfW
xTMcYg+s5NiT3fQaG9YIEQJXF0s5RGMdMrgoDpVs5+PJZEJFNE/HFdpwq12TdhliVAWR0AHJ/EQl
nGdfs6YfafIGGS2SF58MewHY5FPLOHQYJr/2CjgW2gVMrJKgANzRBA0M/30oPeiWMvLMcblnTTNF
LsM3Cg05ICHNimgegyuujAIDsfzHUybuBakj855IDk/p6MkY8z/nERnpmDEebZAM1Up/rsbgXb9j
qowgqs8ChY5yi9Kb2ZSzBlIETJJ1C3/cyyA87kuja12m4mQegTAd+XhQhTUYZgM+37Ns0UaNtA8h
7NtPu6nAp0/OGz4PhmULUPwcZ/TXHvx8VznZhIhdbY7eIZty6LaqDquFPIoZSoUYhGy8s1SWTI8L
/6lPCW/Y0aq3oG2t5WlVIrBtqK59Nw0ipun2WsXVSkx3EuAjb/+QENZfvycMR5o/w/kMjIBnwnlb
qACcR425f8YRpp/sUsJbfEgoUfQvOz4vp97oL/6eOlpY6bhfSGxlw5E5go1IARJs7p4lVcqhXMm1
pBC9b2xrnNu5+l/uVd3ri9Dpz6bM45eJ2VccqHiq0A/C+ftDo93x+JVjBsyvKPj5k9qyCicJXQ8u
7unCcGGY54ADBg8VRiD+twmYfgKnIIJFac+Arq6wmdjwbhZN9HrP0aSFGpziBiq4T5O64PzOERwI
6qFwVmP5kyB+tpxxnC0r/24wZGS/6gF1hR0yNyYOcXt0MD7YZqmtDdqdEmnGmJDiBOnsHVyermoS
8GnyCMYYpIJahp+qWRMlp8NbluM6lOrBCLNKyZZibFoO8KOgEw7GSTebE8UAv84UNVz+PDGeySun
dGtdxiTe0IcBz883dL42O6SUroCN+0yalr5iUjOnbFiRfhij1o7O+DQrrpd7DeL4oWsTV96cGGWQ
hAd2i/sXhygyCd8jPGZMb3NksoKDt5PL0pZTjl3OOX17Scj0LOAA4YvYT2um/4zAiLBn1kvGy0a4
wAhGcfh+3RfiWe62xeWwtGJMoNzMYF7g33NO++o4i8WKug6cQweXd0ND3feQF1/AvjPPrgzmCUZM
6fd8polYp0yTINvQH91fqTXHkl3dNowTtbTxqdfRt6rQZ9QF9ViUAVCFzQx6fRrIq9JcECu2kVPv
ntpsCBU54joTXxm6sUdo/KwyH5byPl6hLnjLHS6LKx7/b++Z/qLUDSDwIb8GKzXnN1PKS6FzQ7dF
IVdw/9G6vBwQZwwrL4lSWIToI73S6yD2Jsy/HbxbnyLAcym6CVAf5ReDsZvuoktYSuTCoKRUFBPH
BhNhUoCm0ZKAwZYpg3XYHvmntl4JYIYvS+2kUr6zVigeEbtdWzzieTkyTWSlsbFnHK8q/cITiVKS
yulsOe8oWWKnk87efeU7v2ShAlr7fCg2VeoLaKEa7msirsd8G0FtMX08p7W1+EDWtT4xPwaEwjmC
A3/mFoERSw1s5NYpeW4yArP4d2c3T7DuDnWl38fV1Tieu7T/i4Iar3eznNCiABXtg2HwGU5cQxBF
Km6S0WVezWb/ujW8t5vTpASEnxwneidz71DeT2cDGKj0xibWQ4Pbk9CkG7XB9sP0tON0P+e9OC2W
oiHbfjv5pDT59Clxqc56z9AiU7AUlg9GfJ9GLfuD4LLKo8t8AfwO+PemNj6X37zfa8TcSKL5ugtG
KXxKaCNIpij+jrKEcxuQyHTh/RCDLfOQa2VaZtIyK3cZjwQfU9miuk0/fh7T/4W03j9OATu9TGJ1
gbuC5p4GawOkC89iQWAVxuWJ0b1kIcPj1GOTz9/ZApI0ZPX19L7Si0dUQQF3v7UltrC8BU+8Govk
Y6hwPbhGaYr8c7WzyQsUHfdFAH05bS2rHhB+EAjaHzeBoV2NwwM3OTNqkPYH9HfIr1dMRhEqukgN
kxe55Xccdn4ebttYydyYPoF0goFQwbsPBnv/I2ib3LWQSyLvNPaYS31icbIWqTH1x8bNNyqDKvTB
0mzAhzLFzawzT3+qyk5wihRzgl5PQJ+GlWb8v43u2CLdLpl0xaElL9MXobvDL/oDK5022RBqiqcU
6dZHRPmm2TuAa1MDzZ1QGXOiqhO+1L+JP8Y1NBR0wuaan3XDjtF9pYgPiyDC48Bv3BkDceCLPzTt
bDHVSaxYhhYNtpX+VRF6XmJcTZm+xBbYHqt97BwKCzOWqW7LvD0ReRq37NlMKwq/H8NZp6BmlNI+
Utc7hHgNG6TVfzV2ObLU95MgRxavJ7fRN4y01YPu+3vZet+zUg5mOgF6Rlr+lrnSfk1I8UfQpy6n
Mr95Ue16Nx511JjNJjoStIUHoTuLuBvUNFq6C4BKRQC8yaXiSfICxWkOjqP4a9uT96Let07h4uX+
hGS8zNnaEWfqcKuBJ89ga+00E13dGLf8qZ2I5pC25zwiBW8ynNjjERkXiXnKkYEMUF+u64HJLCyw
mVeV+gqg+xDupWMqZLXJYsr5DLIx4uniV9nVhcfrlxd4zzROx0sN6qtH4/dBR9rR1nuc6qPd6eEc
KVUAXHeRCMl4R+AxPT3tO05Jc6nj4X6T5JQ5KwSkM0I1AV7skCLXnzxk7n1otoYOS3ZZyddzuFhX
vE/K1pGhOFg3pI9oq/S3upfvu0RD8031wXqm4U42d2kP0EC5hJZtDTD8R6AeCzg27PrazxLDe4HE
SPBKAoI4g7wwnafr2ygNK6mA+oFGpMI7/WXtoShaKIuMN6BFfCcvCPbIQTi4Z0exq/e3lKl3iLa3
euUCbCjncXqYNVyX0KEJ2zrIamei1kS8Nh23tB6woP9R94Q4wnfcAvmWOS+RDFhXLn6WawF+hR0N
tlk6jSRG8VRmos6KrtA47TTPj0mkfDBBTD9+cNXnb1CFGhdi2FZSy04LMrAqtwcFB6woYQPd0qoy
REX5BqvX6VgszU1xYuRX9DdhcsBZOudT4OwuVC619HXkuWuayl/+abgSc28umpSTZU4RaDMBMPig
H1YPA98Lx8YVXoM21ctKd3usyV+ynoFTBl03wqxtDytjZBgJg4qsKram+ZhS9CMGxlvi4xeuznhc
RO2g2GquplTUWDuLjpFUOnv448fB6UHdvCpId1O1hkfn9GmTZDK5RxWKFF8drWh8OgafP41GTa+7
fBSlfWue5K9JWmwLVZ+8OeawuRpvLlXdRDPo8TcUzWwETCdTvo+nJcSeASWnepD2P/n3+U+rwC+A
svczLJjVpHiKrpAHipvXs9LKvAHc/2gSPOO8GB9EoReqcH+LCV9RkKSjbgbKeDfY+Jud010YCAQW
GRkK7f2vjPRsDL7B6Hjm3/BMqpQ26TFQIJ9ixMCgAPOUkONJzJsOVgKNJSp65Z1vW/vEkx2EF3cD
6KRH1nZHpDJ++uWXzm/dPZQd4e7LXeAYFnEQOMp3LzxGXdHcaFUaiiY1naD+bx4IiE5cHZJ5E6iD
p2n4o63djeTTsCVfO3CTUoyqBQ9S1qWXRe5GHwCJloTJYV6U8NS6V778Goj14rv8ssOPgONzhSY+
BWMLsOghOh4ijwDMrurNO/1ZysfNLZROrCTrZz0X40hgw5vWVzdgauUEN8fmRJySxNiSXbL/ck93
OLctCuclrIGFoUJ5GVTcymB/oXofKVkWjEyaWs+dp5tDPRcVLuNaVn0L2yz2cEe73oJZZ8W0E1bZ
V2w2xV56DmSg3Ke8l+JdckNwxyfXgzjesE1Dgyy7L+9IF87XBqeQziVmPVWp7muNNM20zekcixRs
Va+/C4RVL3Vbzu3FNvpSt0eZVL80qoJWb6v/XLchDn3U3I9hcnqnJLzqorG9KfweVw7Jc3cRoD2F
XSH9S7Yag3u9tO5QPVGdjCB61f97uSH/gYdSsaw+8bdvRF2IcI2Pgq9umJXIFHGlQEkMrq8orH39
MDVoZ/drjr8mYS4XNiW+k+bWHNwbhbcN/7+8w5T4z9VEARyoTAkNG2qn/kw60lqkR6rfuV0Zs+ZJ
futsoFIqiQKNCvCmxgqKAldUtOeuYraUkORn5qciNMnsgE9l7aX2hVtzvFUAKe42/PmoVmE2wjED
lN+NqiiTFhY037OIVrfeaWBecR2TkVk1WQSR1ZEcgdaWYhB1e99xx89MlsJvjQ7NKCK8E7cwJ7nu
nFaNkzh8GuTkGJVSo0CnxK0xhJUdHc5wSFbgPBWdBQcizWOHgVPrLBxZ8JWdP2lARxbnQudokEFL
Ca9pj+o049C0qa/9ft227siIeH+fca331gno/1rzAxfvZgQTlgvNfRyhq3u3V+pLLnWbvaW6Ny80
j+xlXFFRETlsXURHxyMYIgwObWmIfGs1brKhgYV4MfsTaV5y1wReh//wJYseSITcTJwYPl9ILRA2
P54BoS8AivdVTjfbMY2ZLm+VcNw69ACLyeQBvjmdt4kEx0nMIHYoLqgdrGduNG1GMsxo8q6Z4+x+
JTZaOEVYFpNjWpnfQJiWcEW+Nf8oLaXbjwUpzVePwiV54Qv7G4WhlyDvXqsBmWN7UYKotbb5rTSY
NFapBmLaZwngLAUQQH8O+pm01qhNJiVklMVrDSE6rSPHjicO7rDAharSKuHJlmNnVqt0gwT6t0fr
/FRgiUyTHrHYHDUlxJJlfY+0yK16wkaDvKSLLrgzevDxqBwEJ0B9/82S84R9nV9IwoDaYP2/6jUv
rdZlM/9FgyfXdQJ3tuRtR8ZUSJB9IChefUdzxmrdR4xGa8CLYBXNL/Lm6xaY1FfNfLp+J9lWl9/m
rkjceFLn3ty/B6/eLBBrpasEy42UeMTn2lEyXBp/s7y2brRKE9PXT7XshvNM2sy1W+RKdUY+2daB
JTbljIkHvYB9za6Q4J1pVtgCBKIyPmbXadLsZFnAEe8gl5JGGmzNW9Nc5mzvzT0uE0H+BOzmy77a
TNT95I9bzk6f9JShxmGTHumt8+mJ9VzwclvNV/UgV9P+CUntGhD4AxN9kaLIUhiE6lJ+1zIgsZ0v
JazJoWrvNXCduKbwuocb6D6DmyJaec0YmRjTiFSn8b2jkbBcmJbPeHom6RLEKSbckFRE+qHbogVO
1OCihBVSObrFKxvztlGYwVh72Z4ItygOZsLEtqSDzCgGdpp5BRBeHDRgHOYg7pXyUiT6Mklahd0q
EDMMrChwYL9V0lGMJqkdDQoe5zyANOHq6vFo+BPdPuCQWOsuvt1TM0FMas5AkXtuq5mv6b75x+aW
e77HqUy6ZCxqPySJlQFC8vw72XlMzddQclAQOc1ZJVDTFujNfuj9UReMZumClKXXx5XMCz8S3tfc
sUHwL62CfuuMkL5gSLkR0/c+uRjH5/4+7DpMRZEPEgKrZnbiAEIxQO2KqWj5UIOy75QNM3xVKQ6b
2DUtbti2BHqBqDN1TTmZ9H3bmvrglKDTKG3gzVTXGpPObTZxdcCZ8PxO1XnjJc+nss1dPzH6oHAv
hhgQ3ilR1sAkqf8HXy5XBY7cxE9GtAMVKKoDvrp2AjzN4MuOb+x4frnL4gjhlgqOH0JoutyOVw1X
aztr0WI3m7AksmzATB1yamMDEWDjDC65KS10AjfqJUjeWQ/HUMuJa4q1GmRGojyweScK6+LjbByd
vORKkF4uc40KhNBSGNkJq3B8CB8u/5H8zzpeLlFPJFpa/SyQ1NeYT51tDF2oSX1ZjiQmYV30Ceue
pxSPGWVtaDLONAfqWvicTxNf4K96cr1ls5iLWy5FzNEFrPietPmkpqgGeul2ql8VwH2IMvSQPJCv
L+e+WdP/1PqUSB1tyHllz30V9jDgcU+2GPTGwWP3TiGUBGko7x1Ja+Y9RFbVNdr2OshkWFPawHO3
9HPtoC7pCtKYWgsOUtp+VM07apGXZ4bJgWPh9q/xajDFlprOmlHndi4fBnriw275Nb4cD0fHZ+x/
0alBdp4tzE/71w8P1ej+82I1++d7ApjjLIzTunicYY2vW7tBYTZmkjAcy0FQZp6g4pz2uNOb/xYJ
c/BZWpfBrfkLQVHAo9jKTypAChmP5J+afihX2GLYcTTH3miJcSYHGFgNu9QOFI/9MQ8rOnZRPAkW
y9X7qrn62KJbRCiFPa6ICiMucUziYczqeuZZtOh7jMNs7FCBOzM2OoEIbtTlaS5afKg0h0UYOenk
qDAppRjsZocVM9/q2xLGwlw53zKyHcRho39v6brFPsX+JRmT+ZxtGndks4F0LSmIKHyc09+vhR0P
nIazx4egjTg70nlaQ1fzAvOCFzTUuZruykpS3RxWPVj3Bvq2Ril7wilk1fcp6FcOcxqlNJzSKgga
w9OQVEQ6xr+G3sTokm82p4P23TyCHK1dNObGn3LXg6Ep7qHjzrl5eVs8VtmmyWOUjPLGRP3k5Ny/
h1joDgFFz0+2gIly0hJOMgFZqXh+QQdkpKBLUHwldcm0hjfMYDls3bv2NlBn7shuy6agHH9wXbee
gyspTCYlK+6PKMRXGtsioR1nv+cLWgrcupSI31HXd1grKLOqjT2VGLtNe0N8IxdFu+K9x6FxAhC7
JSMjYri4iz6oWeQSIiVLNysLjQ0f9aP9tNOxyB9IM8psI9CZkXxsXGaNpdvgOqQcmovGIZasPKOO
DwC1ZEIuaT2XWQc411zBGJX/XdFglPUbtlJs/hvw9+hOGakF6v6R3Q3D6dlVEGs0TUNLbKsw9icW
qV+vQn2E/0LNZcIm/O1JwncmfZWvUIpVPLV4l/FLpOzwaPaoGAUo5ygKHS2HmQr7UZfzXMbYbzmk
WQK+GrWD267ywXBgXVjfaCrXDXGfvZb0gq/CmWl1hjWDfpPZJG5yQZ+7fs/qym4BzU86jITtbPda
fW6VYaRVN1HlML3JZAB9M37hQiVd7FxKWatnTyWATjRVFUgFbepP8G8lJ4J51wycx6Rji73ugJDZ
pKs7bMGwSYAa1ChcIIqjl48arvs1+8ORuDSBhP7TUhnOYFcMsF90DR65tFc0YxDpMIT43bo/4mVD
Y19p0TroeIp3Wak09Bbk7TL4GY4pENV+DGU0X8Uc0HeogjQ2anlNtJZSi0/59OedD0KAG3X973Ha
hmqfgy+ALyw3HNThK5FTDG1bAoRyp7mQdbuM2cvubKEbTIh69FaA6HkE5YmAJimG4HDGqiOdJrkd
fOoS4cz63FWZSDlp4mDr1MlwP2wAc9TwfotP6dfwHChiVGhS54Q/SASdex585q0UZTRLW/FRLYBI
cpI43Dy+4gqaZ+MhZFw+zMXv8hRSdzHsSaGVVrYSArGoUWCGZjsQLTSrJpga72jjGRaQXXx8/NdS
EWBiRLJerJl11NevGvPQTsJpe9KbCZLjTbk9KdehFOHCmzhi8Tyr4gL3V69H0uE83LCT4nBSPBjr
y9cmOIqVcJdluTyjdP61Btmk1d63eFkUICLEBRHZ2HUZblxEoHkdSxHONsNU0fV/M9AmQXzTo+qS
44hNASveTVBxF73Vl6x2nban7VLoe9Mx0+QhIvDYFc9jkg/RYERvbwP/LAy8/wBBVXWdgdKDZqSy
QMx81XkvgKnmoFhnOPyBdDfOpS1KKLnyIEG9l4sZrq3os5wXSBZgMP1AuA9+qbFxFmVDfRXuhpBA
vf/8w88y0W2gQors7Kk6HcfmMASGqtxPAcwsCir6loHgAcAkVAttmvcP7iPyxYoHCR5aU+yPqCU1
/HY36T/8zt3ze2bDpZq6tWnVbkhpsw+IDsSNx9cyUjCPoRjGugXC4LpZ5apUJDMFcNmyxrO8/JsG
aJFI7vQyD+vn+J54V/MhPOLvUs3pVvPthkd3R6KVlQyZzG8ygpsRl7ejc/zBhZtOJtg6AnhSDR1Z
oR3gL6WKk5F8ZBYGEUTs14DugYzDMNC8O1XZ7fsm9W9P9IFb0LOixzk2YZ/qqpULKJTkcaQC/aOp
eczcTN8uM+hepkAPob77lwHXj8bkqYWcgsHHai+UXBlPKkmdU1Zgpd0Sm7YBcihgQ2yyMXgaHTvN
ax3enNZM8LUvFNzLZ/Z7dIvJB3hFtFNqgecVa0xFCVGCNVrd4OXQM8nZ8iZEX4s1IT26A5MVgcXz
NL6G505wSENwWV9UVFWjSPAEQGIBBNOqsaSNt3BnIe2DWY7BWMgqdsmaFfQaduQ0RYhL10nkINMp
TGj03kB55CDNm5ljOmoPCEZWXHy3B9kBx12+UcU3OzzR1ZYG9/XitZaJsJfNFvsqwcDsDbavWcaL
cuzLl8ubwGrQRYPVQrvUlPD3nUxhiCG3lsAfmv++9hkq7rx14/zxSzNAAbCYqxqww0sAX1B31Gje
LcpZ7g10s7/Va6H8wEJV3t5/HYPWLGkp47RqwBjPULByKTcYCsrcPufE6wbeL/UAiqMSwGGWwh/b
8aPGqibB1Dd3YM9ZOYf58lqlxYrWg0wqiS4saD4i7mk2L8dvh5/vFOxDdxc0/dzOxIxScrJDTXfK
+8GHXYgj4WynUq/Nt10yGvVWJhdkplTDVbzDhAW3ok0Y7lH/pH5k7u3uNLXt156fnSHlo7raekpL
wA8u9RTC8tWMzt8O9TFOpOILlObvtEfdP7Ab+y1NEmE6Gu+tJ2g2G8Gmb7CpkEOMQNZAHMYMBFFG
wKKEtz+pB58hie6bfHu/SzvBp25huzOXA2vqcyADB1vtcPQKtFEm13Ncs2geYUbXZ3ABGEnfqn4I
1W1i5iqJFfvZlW0Z8VyjI3DKQz3S2gnBwQr27nS2UFQzyOh5H/2vx1SAsuZX1pkYNBMxctgzO/Lc
OaSfpEYP+bIBtgquLdIDwcLRlcFAuaCnAH0Am2dpuQjH3CUKyQ5j/IL5StlTEkNuJbWpg8UEpDM0
QN2MCdAnaBQ5jtm24G/yreR7ZKDamKzM/4oUIw+Ly0qYnpVZ6LCN45tUA8BbMepuq6vDlaboKCl6
dSqjyWJK7Di6Ok40cox96Jh+6matjNcncYh50O8TZ+972D/v12wpgcy5uk+0gxytdUva9TdgwGQD
MLGGmqQZ47XKGuUVIG2A5NOhsfsr3Ovedm0KG9lEq+lFSWE23i5fU36jO8LPJ/8XRBoWK3iOfDfI
jLVw8TgD4C1m7e/6KlPKKt1HFeh5Ktwn5ezXLlsyAxRiDdL+rbsmR4oJRRZbexfcEzvZ6wVlj25T
4AN0sOf8a5cwGV4BnDOLaDLvgwJr3SDk6fDNloTnx2+1n+zVk35xRRrooT3RsEgY8+VCdvWVf4hy
p8EmcACpVtDdY9UmPaVVMeEQ7NNvzs3hI/x93DI9GzXT+fjmynjjO8lL1fQ4WNwUpg08T+O7USZD
hM6oaqEEipctVJmFJPIKKXYyOgr9lO3wmcIf55P5dmmVFs8E0O9xTeAY6p3yH2Yt/FtBqpIOfKrT
Mg0Jy7DGfNVp2xEp3+aAy2EnH6yNWQe4np6paCdsvdEVUvGRURQ+f8rF+dKW0THh5jPR2rn6mrjp
ubxzMsUlu2elLAx2lXKd4C5R0TSVZEHpVitOG+0WtSz+y7o9Y+PNnYw8a0eEpjW3Ek3s0hbOIeAw
YCOMZc+hXhsoHBcAVfaSqdftMzHlXFsA9iQIOBMgJ4eEI7n5VFiNqNwC9G3gbejF7mleG4qFUq0t
cuzvX7dmpQAwmrwCpG7pc/oIqimctBoprnZMnMWTT6csKOEyOImoRPTFiaFx0FZCTiB1LlhKNRqD
j3Ykbdj0g55yS0CWCW9AwWoLwYQxRkS+/tuT63xxX9jL2W0I/jANj8CLPeHGrmSkm1JTEi2LXiie
C6TIYuTBhQMHTM75qz1jbkR1qRhSqXyAQcsKTh5u6JsHTZQh0CSVXXCpufFsV/ieweh7oxCFAasn
JPuaVjloFCxwUtZukYIHXAJceFms0PKrJckNQQ8/8lQ0J4zd91u5adVKyTqPUzAdosxxhZ8lLRoB
pWm2eDDOzQ4NlTJFs6aT0d0ow7gJgnnnyBEvAFXY6aSIahPyXifa4e4k+hO/jF2luDefoe04Vk4Y
JpqzOK0RjySFFSx8IcB3RrZCePOhYlh2dGwMhRGweLeJnSYv9wXwtdecjhSj7/k7+BdgsDtNuEyP
KyEhancMuCglH0txVd8oNjeqIrystZS/vYmr1b/m+bdjQuXdNrvk+DHrO36MIISBOxzcrnA2EZsN
nIYCujwr9K8f/7shBVAVqAAv8PSN8GLdYss/bWCij08u0t8tYNzSa8bhqSSV+Td5xwdPyS8nWHJC
+EpnkX2MBbBsxpZep9TDKbzA0dXKYXxgyHhWoTcERwmHWVxEq17HkIIPqGNwMvnUPVU3LjG6KHZp
AK65b2eA9C4bQnqQu1eKVSjqdogbpVJWhgztDZFqlPToW2Ctha22IgkvRpEuDw9juprT/kf/eU4Q
gPuZUCLnLAS+FpnOaOduZ+J9ih8RE/phTq3IksWRK5Excr3jPlT6GfdfXuvGTC1DFvQ3RLzFknuN
kqL3t1RSTIMUO+HVgvKNx/FhT9B1aiWrwg5mWtbbYrxzQqCXiMfIJRVYUJWM6NktopOO2dK/JIkV
ztQfiImyzG6HtYHJkOM2H+vhvcQYlLHBqV9RxXtXKxN8/ioZFE9x10zQac4OGUGekxl78bwCHato
1Iud75K2ti0U4j1ymglZVFGEkWQ3+h1I1u6EX0OZy148OMLwcP7K5Osq9jlp+lhMfvT3vYYjPCnM
bEuuZVrN0jev/8ScOru+nFTDmxBEvCJcn96tvWzwdo77fY5616wZgEwhWCrvsPdMQU/GfRj1EJF8
LWgUpUPR5PJPFx5Ku9smulYUUhw4mVDMjp3H+h0F328hQ/JapU+M9IxU4x5iQlPWsUV/p5/TIwCI
r53v/MIbDzzDaHchxOUD8QxoxofsHc217JuNfamse6v1z2AlpdpL+gBQq+B8ouHGLwU4Xps4GTSq
Zk41UcVt14pM9shopMeoxTPd79lL39ltpxMvGuP4FZmVIv1JyLL9qPbBvl9ZjFOmzHbdhkPjGAWg
C0VC+6xwwSs85uMsPZ9LQ9o2WXNgG+Hkl1iWSxbUrXIIvtSiKM08gGYJ+0n+SmDme/J8k6QPD2X8
X5Q918yA2/7GyxMX892ydJy4i3CRZyk0SAw/+FGu8Pmy+zVyqIPKqGQ+avJ5exvq6cAU2b0JeOaL
RByoaoZIK7jCJ3qi/AD78PSPD/yuRh5XCcAHfjm02UZjmhNmdsAHBcKZThvCQ6eXE8WQ1HdUI5Z2
jrXHvlVCIT/xf6QJDonYgOA92+t36xQgX3JhvVBm89tiwiCDVuoOqU3S6Tga79FIHSU2/CmtptIH
/8Ye2Jw3B+boasMC2Eayd7cvDoZUUd3g6pnMKTau/HfPSG+hFdu5CkATWwc11ZpFtc+xRKgEpCl7
ioPchOVzOWZWrQPIYHNtddrlzxE1YY1/A8dBvoeK2YgtrHytHBwwRKEaBQMYrF4uwrPGLQKYFJQe
/4UWpRp/wg+Bp8e/8l58lbadXxtZWhy9SgKMxpckD2SxhT9+gMoPBB24KBC9v12Jq1KaP4MvGgqi
tYjuvL9cbxJCS4lamsC/okNvGelIJTCxFwh20kQNQ7GddkT70LWB9Ge/woPwquIXjD7KEISCs2g+
b82gIoglKZr2QCaZf3QaPBw+jN+p/z1denYaXEpFbiLryAcrtv6nXQ2zuYCeQjn3GXG9LHfl7i+h
/i5+QjQhuldkWAJLtPx4+jIyd2KZjttpaZGhYLhkgVKVImu7JbkJu76/fqadHXcLU2TKJF5XxJUP
TrgehdMe7W68AeoBNl7uacnBGf0vJShvSDxM2H5sqLJtmDCACZ2yDWDYZhiDFx3L6L36bFqITVT2
y/YnoAxMzOixL9O9A67PYcfu/nEwlKKIOn7SNLupiZiQTRfY6QqrSylkA2vQSqLQkCKVpvSERwFj
U9BslGZ9To3vacTbbSRuDVmLwK0el7evsYZQICstLyQLept7xtRejKIFMIStSU74lmFh2MJ78Hon
YpU4Pse3G9q80mPpqR4mtnI/mYwPIsgupnZsQFNHREpAxrFc6LqHbBK/EuSvb6HBZ8oslWYeG+3j
Vc+HXrKWM4sR0Y06l83bBeQs7NxMFbuI4lnCSUb3uXunu70gI3IWCC0oi1T/pof/t7UdChARsAlP
cN3CwnpYqrCJEDCaUe942sLzVOUeNInUHWo5+qdt8ty9V2NYudILq0jRM5gPxPdNww6jDGddSp3W
w5WqaCr/7ncw54ZhcaOtKkKOAGlnj1JLaFsGXXlHIRyKZ9W6tCNryT6N0jFtHDgs0hAI8tcU6CeX
THSO1tqFpq+JiKqs1Z2Mo4JWXBf7u2a7JVyKy2RaUxWgRGvwDMIZ3losAiFWpoWWI7gq7MbGBUYX
/OUwpjHKR/1dyXsDKkzawCoT2cBN4XLJTnJVtZaWSvkGD1cs4sIueTNwjptd6q6goy35BNs6/2gl
ofI/VoSC7G/B2za+hQhd7UTPLPkkawGf5g9iUg3K+rgguK+NEOa5/mwcYHHhRfhVKrHZ/3hKkyPZ
HMp9lTxEOrsYSX/9WYdfguc7UalaozZtptf6XyWK9kuBgaAZf9aDuyMSPnP/QCGqi5H5tf3y9Arb
eXKAhlFfoAjWZtt+AyAJuyzzThUrtp2X4dZqB3X/5Yx6MC+YhPJCHGBUYOtsgEitxt143gq2gms5
wJqg2b4R5pKrAx3oxcfzRWLEbf6n68vfnWHc1aQQ5LdsmBuuIh/f4YKiU+qcwDV1m3OHcoMc2K7Z
Jfu1ZpTRd7mznYVLO+DAaayUI6bwKeyAck7u3zDTvr2+XCYW7/PhBLs6RZ1R705K03vw4h4mNWx4
tlWGJavyoRWI9WLCi3EEQHJgQL0UtoIyy2uEIFPWXValQhK6bL6qpe0ps2WLztl42VwUQCszqAKW
dr4Luum0376tR33vWQkL+uldtp2sU/L8xpt9RP8V1wm2pJGqTbolZOPnmy86qA+ZmuauOcbeemWe
mYHB961oIywasYswOU52K25OGxqBuO0rutKdU+1OH/ceKic5vZpCX9Hzoss+VqASjK5P1gLlyqln
lnEY8+TyOP1x/qkHKBl4iLjTRt7Ttnia4rVupGGaiXYu6+le/veNFTpHfcdsOm5iDjcYxOVw2K9L
QlqVk31Sx/FDUBggGejvhed9Ylk7cRM1k9e5sfsMedVxo1k3kEkudiiYSqeXNcfJOVU9jRPYxUhe
IzAYNJ1e8/NA4Zke7rccQ3ylFbzK060guuFQcfCK9QkK/6Xet1yP+ONx0J5rwP4L1NJS1Pxr5GXQ
hEXmEaxmiPK0H1+I8xmEhthymDKP2RBrs1raiYZV0chKl4gfyQuHNGLknHkVEnd3BxT7dFxk5RKM
XBv8ABP5yBOec7zPkgYbDjwxTa3/hJZb9UsWqyp38Pjn5qwjvvjC4TQ15OXmgvp65HZ7EIwYudKO
95/HcyIXZzSoag4SYFd0cbblXL9sjCdzlIhPEJlKL9/E6ix0UdxsJew7pEDss2BbblNZ/gseLFxk
SozbfQnO5k9ezd0brZceUjk2pImmpvC5r6xU0pJvOBpb/9Rbd3f5VvSwfR6NXgo2EcC3LGqoIyqk
wWoY2aqXuOqGVwLk5Wj0sLjG8ARbO8iXymMCj5oiVuZaZ6yU9/kXg1YIaBmBFWcBOmG8P1Rvd2yw
C8682i2r+VYMYZVhdPYXAg7RjMbuxBjPjAXalMwyqDq3x5JYelOOlOf8vH6cCfT7fMwXbIOqZJ3E
97QzCQ53jNOie/me5HtvUkDD/m5TIyBQ30Gb8M48av69+OzAhsOPyjOHVGUQQycnQRB0ujbHwe23
sxeB3rv6G9jNo4Bjst9qdCyUs9RhsTiK4HFwRl5Msdad+eoW07dMAdfIR0VY3goUdIoyvgkWanyb
zOZ5rh+OaQAvm2XtzT6PC13MBvp6hX+NiXFD4kAz8x1PtxL0P8gXCO83M9NzvHFr31Relh1wMBmO
zdO9mEkPsh2DyW0+Dbr1SveGmIUgt0nkdjMYKYf/XQgWq5HDDlc72cK0sgXrV+AbAnBRVvrHiZNo
U+G0lDFroP8cJsf1wZlGm7so+ym919YZMKJj2wLDTMxd8MrdHfX05FtWCKMgnwNJHRvHaPy/ngXS
yysP0HXMPPaRT429i4+lVU2ag+GleR+ZGYhrqp30aCuQCtzb9qXLFEFFCwHFHJaTtWOsjbKuax9z
I1HbrMH18cxj9MUjSFrXLK0bLPQaya/isp14W8OcduIVZWU0rhI/5EWV76U62pr1ZK/j+0zRAURa
jf8+qF1QxehYK8GK3I3E9e6EYVoKo4K3oY5n3XPwSimgYvHyXA+vhsG8s/lyF70cGyCS8qWKi11m
v8bvUrjiO0qkIq/ouX7NTtOD5paBWSVUvL6EQ3+1knmHygwh/aS6Hr4PMxz8YxZmrEdvYxAa6Qm8
ssG2TMNTymhGkPgMl54I3DZJ8QczvdZxpJ5FvO4T/jml8tHxsLKI4voPwJ8uP7nwhFhs3N2EnEAY
MSXYGz07GyDODu2EQuiEbXV7rYg0/B0fvCIwWXpF9ICvWUFIjG2HI1atABN4W0qwmeprfyM25FfA
uIJTgsi7bhsDnudxSRdNZEblNamLjXivunHWkI/hygnuvFgK+FggVb1z0MFI2RM/XtAU1cp5uY8+
b553d760K68EWm7+1CgOjRuao6dxzNyvmA0su4q++APsO3MP45EP2KeiX0celcJq7/HYekduFDQh
RYlv4M7e1+pt2DbIWMzxHXf8VyfFJD6vyqVK56oRrWyoJLvWNGmaiApKrClZYOSn/WFoNT2sCgxH
E/pEmqjModstbb/RiJFB5y41SXFHHWItlpaoFEDITjYpWC1EHiTeK5VfnJLM/r+qMBeLn/CScg+G
tHKfd/3e31xCLD0jPRDPXHgLh+ypadb7AdVTDhbnQmuFLrS+PSKi6aP9M9uISc9/J1CtNTIvzuDj
NdqDxytBjDpTJ35CgSHJopAJFEMYPgU7nckxrLopXUQLkIm5kxrGHlmX0vkV8jvyKNlHFlCQAMJb
zGotn2JQdHDDGqBiKYCNEdQABOVUrYZh1/OvXs8BOfSByUw29N55V4+5JVEYwCmx4uJwtNrdwCnR
DYRFE7CtTdn7vYlE+ZgwZls17kHxokXDB7Lrp8QIj/evedJMstzGSAoni5aDfBDe1N39GhfdjUZW
ovX29JH4wZcHjyuQJMZDm7chwxX3IwmMhot5W84WBmM+Bl8Ijm5ZokGR5P2JBzqibE/XS9+S/kt4
4/ihWn8Rh92tf3rsq0WF96wFJ593DLWbVueg03S80yvYZ5W+yeV7GLUVlS79PFbslPmm443c3FBt
kw58V8r4z/ZDoLEZbsF8nZFUqh0Q/Gud3Uz+ZqUgf3NSkxMcIbxVgt2wIzoFDW0urBxY1GIwLu6J
HBdf3oHlOg+nsVXqlLVF37mfhgb4M0PYJLMepxyNY1tV83R2XwGZXFX8UGhk6lA2Q+t89fe2Hlsi
WhGYxWOWXJc7c2MGnN/CDnzuq9cVjAEZsiJR2gy4OBUgfXJa8Td6Cl66WDgt2HqvMeqtlN8DzTkk
SJCqbmklFOABr1ZXPi5405rjZ3PY719V0PTobdregdvThMBMZW0LmFF/OmRmre4EuYq9DSUeTw6Q
iS7XdMLh3SqCrPnBnZAmoM4aFyBYHuROpk3tKciN7RDg/u+Smo6WpYA2tfe9EMamfaebfilANMh8
hYfBYEquK9qhhkdu0XHzvQNpBw9i3qQXoNQYq9TDNBHpNjMudvW5BeuVC5VTBuzJ3yvP0UP7sCZt
9XQ5jJOL9SVA4fA+AvHDveFNgh9973RAb4rHw/B1H4t56MuAywvygKDFbY4H7XHDB65tc9BXkwF6
0vUwrjMPhtkkSfwTP2aD6L1Pz3NUWINAmruVkuDGzNDH0XqZcFOsRyn2cpssS4fdSvQFfty8ok+z
ri9WL6xPCgs+oeZdep8wL76tTeH77T8cZKkyIfUpMQCb/UQ07AX/hPGHi2iaA3Dla2VyWajMSSOx
llPv7tHWVFxGN/hpDMq0HvaZLX3AFJf+SQIBfBCHa51MH2i95ng7eo3OE5qmeYtCho6WZAoTmoYj
9M6yojEzysg91j34KdmgjPLfM62Bj36HgE7r+j9Z6Es2PpCUKVapFzSyAWW8xNOO+p2waFJz3lxa
f2sr9iu/gAoZEn3PUnm8MLSCMIqIVewPtYlMhlMFc2pCSFzwaslI7lyJ14k76D4FyCcgxB1OCPwh
6ScTHou5OFTGDwKmi61cKY1HgqWxPXX7Zgo8VvpCnTAb/W3R6+wksUN6iyrS/2apq7sawksfrWyi
Ev+GzTnXGYtiNSTQjlqFFO25ycpfxrdrJErcM8LBevXyK+0VBFbKcX+Q24VSEMIBkekWe5YQuwLt
GBlSaKzWNqyq0fHiND1ZTj6WdMbekVNEunqQM65Whn57XArtJcHBuF9r8JjPyNu0nrd2Nl7RKonh
IIo0sUHuVdWpxguw2rv8uhb/lUIJAy9Z7lrCUssjE81wkCt4YF6FhSqJgs5CMjSTy6TcXqSa4AQ5
Ev75wxQqdk+wSa6Ln0cIPvdZyKqetFyHvPtgFupLSTB4ZOILJQA1cXW9ODwDe7Wjht+udLaWMfVN
AIubNIeve27hMTMyjQNMifc7Xi1UJYfPy/zZmZ7HBwASpmgsl06A6oG/APzsjgmXesi0+v/Rbbo2
k89UHLYHxu6kO/LW3AB3Vz6/hjKKobk/puoMXwHM9O2kNFBviL1jVZ3ff4iERF/PNf4CHUWPUNwq
wnad7LflE8z+Hj5UJENCAVOalM9kfcdMbNzO1FFNuHBF7bf0FZoqtqVNBrQqJv6Aht6hyXIWyCkG
goWu+NYAeGAT5yhU0WPr13G0ZdIpu3mjvMtOf6fkk6Urax8gbTnypQbEJ/X7uur0sg3WVR+Q0o6p
rHMrbShCOOcoMWjIGgfXobAgnhydwkVE7+vvFL99+C1S5dkAvE3gbKkU+167WT1Lb9wnXDPW0NhF
KQDb95uxX1ZqqiSng9tUilYsSRUGoxlC1942pgAWGt7uusAq+NrhGzUglwzYCfYOOrLY/DATR8ya
P8myb3sJuMQamGMYN7fWD9ReSNZAGpAYUt90yUHBNuR2sDfIf9sKalBq2d1NLltzWtQNmrG72lwv
F5ViAKVC2Xs16Vt8eESh2zqsjRXU4sokCkJWBH+SXPx1BXTGDDQDM+Lh6YO8fu9w/6U4/lok9c8L
CRoCpsjE49qSgtcR4vED1AaDUMFcKpOSX8y1B98izzDFSIzxydDk8Rlt73qIAPpAjYubmfHhp1+p
5T6bmHp36mblQqubkggf7tTEKpIk6jamepHVSEBgUlLM1iTQOD9uYO2fbhaU35QingSUPVt5J8PX
1HBHWkaCMrpAZeolw1kgL3AtnUyy0le/e0PQEgJo4bCyavad1MxogwC2ljlNtXL7k9eMSx3IYbRM
EhYPLwc4jXWuyU1rTpooAud/HQQVZcIsX2Sk2vVDGfRQPZ4EMVXFfImqHqUGZ3nt9UiT/XYzGbpc
Nuw1u8TsbMbq2eM0pX8zK9LCz5KIvt+wrXal7a1zJRv+9lxnxY6eOopfy2A2druUp2t/Lse5k2NR
/tblBVrjhlJ8I7o7CHsaFJBrV+CqVDJ62vX4uWqsxB8LJLQ4dKQ9hefPTqOmNtWH0yZKosro7wiu
34Y7hevQ/QO+AKKvrPuYPicpiAQwUaiAEtjwht0KNj346t1Gm+iEqiM/6LUQMJ78Xs3G3DAq+LR/
OQVrh1N7CynnOdVGIpNQmto7vcf/l+8fzTGIt9Q+2efm+qlrCFL6NIJHSh5hFuXjZ+PFUVuvGIwg
f7/2+QBA1MMRpDfXrz6/h3IHIAAy95iAg2EXSCYIrrJZckK5wqFKA+rVTY099/hW9yLkthXjHK31
KRKZNzDVCkaXTFxZHrp++n0pF01ZCCH7NUhqb/YFWz9CQ9H6okW9xMeSFYCD/KHTbzvj4fwPpZEo
FTjiIl9Hejyi8oYBgCh5GxXiQg4ooNr6g7oBCH0S4/AUFmMxAOuvWaN2nA7MDfnLh1lLzBoLAujC
IY/0/zEKIRKDTK+/QnmWBiCtcbISoGjafQ/wRpWnI+DWUXSr5k1f8eGqTKYFs0OBUWxarPIl9CQ8
i11isdmG40+6dBtj31Tvmd70+PbfI5n8wZOG89KZcLb8oupWI5aWfnyLEhSxlvncIZwp2dbPj79s
RD0zyxn686HkTJVeSHflEDPAESVupA1/PQQk8ynDyZ/D4WiWAB8gcROpJmntxLv/yBI74yGGABsb
ePW60BiQ77TPvOVrOo5lTOrhILwsEzy/yEyMdG4l3qtaynOrfJHynQB+sSTfWbbwjhWzrDp2Vfxx
3TNPwVM0gDfno6IcqoRLYViNofg5uIyOLK28p36qygcYUoRdgbGfjSpYfX9kJPWISgS9Ce0728oh
KhF2SgZnhzmZGS4H003UG6I/0uR+NnTtjtskCYNSSOu1yYkammpXFwgnO4z1qYWHE6FTFU3HFMMd
AAQHFTsfPuQiCow/6FwFNL0brH9lEFVtMgEiax4PiqODiqNOMyIweCfi0y27bVTLs7b24RQACdAL
Ulmm3ktBQ2LDjwuW7FGonLfRJLjfRncTcr9LQUjkMsjSgAOx//8lct1wc4+MA6hMezK6cNjiNagl
auDpztMReWgC7j1/sQKT8wJGfV9FzRtRE8aHRL5UpV8Eb9bjJo090jmCSpqA6d5dDrbTy3zgWZ4H
tZzXhdDIT3sfCreOS/Hzbu5PWzcOkICc6v45ioxVnpE2Q5oIuiFE4Js3lcyWsUZdhBxQ1vqPDlmg
cFUgtdo3KK0de4RLeCUebHsRJvzXIpMaDMlplUK+/Q4pZZ3Hlutn28fJw4C8JqlkBrjFW/GNQBOr
e9RLQoJZTVN0WgVWUy1TVqBM80X/nw4Ma7I/akVA1W8P98gvTy4ZAvjbobt7DWib7tToS+FmlMWA
e9AaSwJhyHDo1b/Dm3xu/CNgroTfAd+gYfZqjqXZ5J+x1JHzjY/D1zJLnsXorqGgLCAymDEee+b6
d02v4SxCEzfwzG5U1h6+F2MfqqE9cz80aWBwn0JiBdSHJ5U4Xn5tAUW9jskzAM/Us/7p7pwxMKjp
/HUGFv1qDPeFQHnXzYYybSgMZH6qOMwH/3rtixvNfNIn/RYaDO4846lSC0AZDmgCFSfSGTQESzFF
sbBp0agRNQc3AxMp4OFWIHXNjGfOvRhMPFBdHV7mK1S7UYQ0C0fqgLD/sFL1RQ/4aDdlb43AsZdz
tjOWzsTNSemaguMsQLQuaYuLzV5/2rPKYZOCbvb9yD4KkQ9jKJN89miM6CqS0GF9CDgPZIz9bRYX
v7+5AMdL7VcVm91HRWPERbm9dkCCDto0zI6/w9Fx981hoSm8sOt2zFNlEI8vV2dcbRhxx4LdgTCc
XD3EMN2rj1P8Litu/HHpaJZUVfLkMDkgIkmyAK8eCpBC6H47fe7sWTA2xdZ9UMSUU2N8wtn44+z6
zubdzecSckIzvBpVVWj2jeLzNnsuRCNelDk4Bls4CgxR+bWxUVcor200ggc+5QhDtCRCifVAMKjr
RgjBY3JuK9CrytFmcgDUmIq1UrzkLIxYxtOHLjqKkYiofAj9rFLAXzqh7LDfuF1IOcjZBBrHHrJz
91TPOBth9cBojNP1Av5KAzvtohpGnRO89TsrSILYjz531U8V8+X6P+8O+qRb7yFdeadupVReP4U5
MCMRMVBCL93+L8/oUdMnFzGKxVuhdFO1JSK1NcVPAoL9nqbw+8OlLFZOROTvQPOz/yfr3giSJG2s
Wqp1IURzF79uRItjBZI5bg1d1wBZ1YILNsBO0dZFacEsWmwARs6Fenl7+3mm4KsURR7QQJ3LW2CU
vhaboA7/I/PU1RY5Fthhl1eUAQOEf170+dS2cBoYUtYar3Wq/jDH1RuV/hQiHsM9ndiPGpnYx73M
6gJvBIMKcH8iUXq3s1Lk55xJ39Omz0gBnQwwCim99dc+t1FTvsfFV7w83SQxGyM4s0eC1TkJ55VE
6brY5go/RLowpi5JBb4vSQeRGro8nk3liJ/vOssQXbInREjgmS9fbNW0tiIhm8mlAsOhITeQHno9
LkqnoiPZquJqwaxkU3V2LfwwxvqHkmBOD+0sGRvl6JmY14977mA/YrDbnQG/7tCxwyFWj2wr7WYr
BLa8E3K1W6nU8LfGB17buP3+65PtahFdnEcoOuQnj6exa305cMsCQafSooXWH8BqFfAmsh299kaV
3Qpvd8FQxA+VWtM5+6WYp9SKAee1Yh/zC+2FQL2fwDHjZ8NO9YxqqZpafhfSkJ8Bep3/wHMIp7UN
YueOP8lJ0ZJ5VtxUTf2OXZbNv6Qu4YiA+hj9UidvRZ0enQRzsZ/9ODC/TkeX0X71rjwQIflRWRaQ
h9qdKcF+9kYo5chpuDHqiZpH2NmdobmOf39hFTv8phuK6K0IfghibUZMAuv7bUhU2RIBfrq8cOY/
Ef+6F4OifV6WOuFvlURfHO+A1GWEatDYVD+syq8tWLz2lbZO0Qx4aPYGmJkUv9ZvPsSH+AM9nirm
4+mWVKNo9BrgrVkJMzhMpERz9ChP/sWHwhCvwWbDY2F/SSRraBlx8RtmJNQ03Ycp11aohgsMAtHk
ptXUQHaddGwVNXjHsfo6HcTV9sTjw5I+t0TOuBjVHD9PlI9T8ci7189s4EM4+XxWMxwmIJ0UD4wb
fhcxdhrJqHeqBPTY3a0TzPg+x8KKD4fzbE+l0Nmitje1pbSI4Hcs2EkNUsb+du0QpFdwaEsCg8ph
s9nzRQ22Q0V2Ai8NmuHuqrEz0fp94LEYK58uRPgizq2uIc0rNUYNRKQBI2WpEu0b1hK5lehEd/KE
P2XhidUiD7bPYpYsBgwsvWmwvC0Mdp8dj8pvSqLAsjEfpEauORS0u3UjWrGVbz/fabO4eq+vGmzf
ufYvkBlrThqEwsNGH0Gnpd06QQZ/wzS5quwApWPb9cMrVbpF7sUUuvrSLUJVz/kxMenTX2aNynub
MWXGz2HwCsMLnVsV3vypdaQ06l4ngpAFxGGh2RJAZgXXnEpH6/KTb3gQWjR0Nxeb7lGmv3VcAnW/
9NlqTBz1qJVXbKeoXdW0oYABCAdTMu/zRys1rt8vy9jLnWtbjzNBc74grUsSfhG8yQad8hR6HPGE
yDzk1QTGEe6me8NfEIBh62xMyz4kS+wvddB+kz71M5qLdtO/yEFsLRerY9dYBTLQUb750odeP8LQ
LcdpSDGiarGovlxYbY4K/KcAlugCvqsSTvwColBusf7NEB+VXiLU9SfD8PONiNo/ik0YMFUgZyBy
dLADHY4AwwawL9kZ0QxjnixM+dl9GMTqzXJUPqbuIygo88Ls3qPIrUBgeWmu34/bwbuV0OvXymwr
k2kNxKq9NMMCyFze3lxKxvHkyF0zmPrQxJ7ravHHVSttd1IfNgVbffx6vdPERAwwgf+XI4jvYfQx
0TVLa07ZNdo5bsxHHfWuOxO73YhGqDhxLcfXe/2/tH7IRBVnN4wy4OW+L5iJCGxEC1C+AoVaFH+u
5e9ys2DdVM7V8pcq32XUDckuazjHcGJRS2UIF0KRh6q4P/75ZAAVmgvDBophdhg+z9hoc1b9vy65
zjgc6JcJObVw9GE9qXdZz5dURyhSmPneAQViUuabo4lmN5h1OlAHJkX6TOimydp2FvjOV3x/50x3
lN7HTRdt7VmUbA/bXhat2GY7XzYfYLDqxjK241ojVy1iGuY9jkJMvKgOV8OiEbP6ApAjaasGDOyy
lTHoMvDHgENu1dLbrFU7txpU7FwWFTiUbJ/WYXYT723Qued/wnB58A31HQFwTdH99csXHcpy2aac
TI8Gguj/Bg4uvazOk12/6ED0sw+SXuWJZeL8V1I1anf3ZrP75Cd7Pyc68GgpZDXUcmi3/pkMvs//
o2CmLggD1gcSmp69VMknE1jWO4c+xOM9oTKL1chzsAz2nH1GivQokgCfvmSFHYk4SyFT8pFukYyz
QydqaPQX9cImg5h4DVJRtPhKm/hRGIne3SBUUq77ud5kM4EicNee3GkbG4muC84fqTWsUs57hIEZ
EjGu5VQ6glpEaT4n3Xgx13nXrQfFzUAPF9Y2JrXc4wPNxshYiENdwq/2x5WGzzEBBNaugRKERpZK
4yjqBWnf5o68iLBP7TCoEcFMiEb7n3KtfCc4sYcS2RcfGAqICPgmWVYPoFXUSJmioH6NYvyrgIBJ
TBwrgmIqKWpR6e32ER7Awag2c/uNZoJLfJSaNQBccdFw2NHN/spJPFfgG6Hi4KyKMTmwfoZy9YdC
Zz0obuppoph4KCiNY8uju8JRBrqnWvUJ4Y4fKSc0avFy1we2DpKjRwAywRT+rupLwEA6MBSaMgRt
FPxA3oJP42RxeQ+z3UbfWFq69cM8JkV/ITqUcXLH1KOeGDZHBDLLHSoRmudrUI/ePBdMEPd+bCM1
/SxREJCVwii0ggVAiMVhRHBRPUKs+gAguSDictftPSifBDoRkYQlJHNt8Y3a1JWq+3jNgbo1hhkD
sONvJyFlgCX5wllNjN4dG3r9W14Q4Os+nAwS/nAoxpljjo2ADU9H0W4FBwsrtdLVh4m6G093OWUy
0SxnSL4/gJH1aCn1g5qVXgvraqzXjgs2X5BezM5nft4Ic1YwzJigRFlrEiP8toysQIuD2R+x04i5
Q6SInVh9k/Or0FhlmUiTajO2OO+wTWJE3pXkzbQqQZyGJEMhzQ6qR/qz1Xl5Jxm3A5r5fSmD8FTN
RgmCCGI4/2MJxeCgt+Au+gfrlq1bJWarUeoQ/q1ge0SHKe0DeZ4qAP0HbCEknR8zncEEHdnu9Ukw
cRDTbUERjLrx6V1cWeVBq8/INmdYNb+dWXluloiqkzQ5CvFrdmtH7vgXkK09ph4hJvmQNXE9ASCl
6s2+9wpQo1yIW1/M5osUFRrs73kOxHuGf7744v3uEYTVWYdy4y9rbgiPSztG8NeI8DXcjahvAcjJ
QqpC3CNqI0budOlHlB7Bb3W4sbbkcT9w1BNPEFD+Ej7NDRJ2RXItCFfpJdLaDRHAnw2xDv8OD9Ek
ZWJim+XnXpkNoWNxCCg8g0FoaKbOXchxp3FE8nonxiMztIJS7aqJw4eYYI1Ma4lfJPHUeBpb9wRZ
v6VeW75a6Ufj77Luhtk5IIy/ChDM9NlEqllxViTW03WePQkd21TSbYyWOgMTyUh00NkVaCZ9h8GM
6gwpFtgJeLGH4plxiZiD5mG3N6alZLjbRkMoYOceVDPwrjh9vz2CEQRCquMK5kKH+OhzmJNNlk78
xlzT3tPeOLkCdDslz0jwUk1vYDEL4nVHqCitku1CcBmTor0ppAD7xGaMlIop9vG3+GsuRwK+wlC3
FWRDaXCv9Cym5vqPPk9gD8ue3wkRyoehOi9PgJt/vT3lZH253Kzwui4z1gu9yB3B6Vv4x+IV+BEL
UiN/gtFYpnp5i5uPHCxV/7vXNAoD8vI+pyONyrcF0/Bh2Lc+brHDFeNXhA/vcIcQGNROhmJ34jbY
Lm5KWqO7NM9CpR4orC/VqwWXtkqP626v38KCEaaIeI9BDXaUUgM+nzoIYLaWNO+DSM/NwjuwN58E
OSn93vUYa5yVONrC/zRXF+Is3Ze/ZsqUKDeamLMf1oruTAq5EKRc8eg/IRUiluiQubqd14cEhSBi
HKYp+y4Z5TBWxdn8q2DSiO3FzbKPyIWQVfepPNW0UWNDJtNY+nDuxtrC7sv2jK7R22tKpGsf5W30
IwqfTmOudgAK9EFhod9GuXDuzDqvvl+3p3/06dtTWRO3I01m2aFRDHZycOOhZ8lYnveOMA0JDHGC
clA/jCiq37zdzEhgDlVxHFUpZ9SXwpQvAy9GLY6ndjxBLwFH9hSmiTvR2FihZSCWJmz9+urgpKRe
CZWbFSlR8ZZuPxr14Fj4i8gdSMTKF+ZPX/cAth8WjViNIVTcYU5S6xEHbBY+NskNUx05W+AFE9dY
djqcc3doNfLtS8JirUZCt54iz3LuYDvJEiAOkAdXVZve5wy/ZoIQzGmlJjehsCkTCbASqsr6XE0T
7UAHpjkmCfIZEXJK7ZJTG4HzQp1bGT7sN+j+trwzA0SYSU0XgDfSzYd+w2pE2Jpp6w77rj17AQQ/
cW/X+NMRWJdJmvJILiWElj2LH90/aTJAEeHz4oCrwWXc++Wjsw4fkn7h3V22D7K2RUBGvsRp7XD2
LmmjAf1tL9d3VyxfMtQZFC/7W2KjJ+XMqLiZ8DQw0feIxtATYLj6JOaGe8gvRRjSMSm13QEjtZuV
7MIsaOnYQ2ZI1UU1f5dikoJYtdxzOOQBi8S8dZgNia2QAfvt7QMIXXVKOyfAUbqcoTggHGnIwhj8
4/glhsHknAeEO2KvzoE9KvOGqTQJTCPWTiWZBvAj3WuYV6KUu5n1roCI4QrJ0U4+YC5KgI6m2/ej
yt6xPKHh1JhKKWYi4dIPEsgU4tmhoFUT9Tz/ccNPL2mdaua+VeFDmh9pMGAYbXePIPh3eSG3R7eq
uvMJ7at/8soAEyFZNLkC7vdXN/K7F0S/klNk1QgSU+Age74SHRHUuVpRrjq/RbZhoYq0IYFduWMN
J0cqqwWMea/T2LR+MUJWFudj8RLZHXRRKhjeLFZBTv4x5qyoZcp/0Uek1bZdMyzTzIjNZEu42/56
9pyfFoXo7EY7OoVANmISCyj7JEUGrlLAaxMmuunzch9ms41Zkmmwi8AvKnae9acOk7zikrrZAyrD
inOhjte/DjOZxEFHqq5Pqe6LDCzE3mpZc6OqgHRL9MaFgP8luEdhTXvlHPzAJQf6gcM6G6gEppRk
5N2SRxmVhlUvIQA7gI1XbNfPGBtpPQScSrFfdgkT6rtCPPxa48uXTQTxywlRZbVLAt7cBVFAnfmL
xwx1zWk/mdO+h6KsVQrvutvH14cf76eyqmoWAuLDK9j7TvPZya975770Jea+PNs/HbC0FjoVanpz
UPoAkjNuMsmDEqAX6HtmmhxhEMUd382ozYvEKTLR3kLjYg6wZoUQAnc3nPGT6wDYAEKPhqOVzBQs
TljP5bIGT7mGFDI6ie6kGk7DmAm3guv+7BWCcl3Q3JaBGAYwSQkD7wYz8vRA/HzP4nGzGEBIKxxF
ZtJ6Zgip5qk66NjY17rbnLTjsE65B3mWM8W0Zax7qQ5/twYqUgEhWIUnvDpUiPvfcaFP52RUWBSf
t0lbsU2mwj20MWXAVWP4QHR5OxLFe5w1JYV9heDhMxHNUQc2wFiIdQv7A/3uKgwF+8uC9HvfJJTU
hFoyhsYRdxord6dndkYIHrIrEge4OtT8/kBFYSxshYPeuFAa9tVdcyzpA31mVZPEZVpQaWvG8lZu
b/Y/Ar8OUOM0ieKArtDIKytNcPVRvXXljNsh9X2akd3d6GTJLuLkEBM47XiX+47oGvKcDJZ9B4iC
x9nKBZXbzkuw+cQTRTWxNp6OSAlE8QYwET4Cl1HIMhpyKfx8IzfGxsnRdZs2srvJexhN8PQ1h/iz
q7D8pUYCkEW9/+4pu0MI6lzKtUCoWBUgGi/AxtZNEI9UDMRTWYO6ejZq9Di6u2a1uc2GL0L+ha0r
WNwFvVZg9fqyqLmpqGNLN/8jHrUlY1QMff7fOvzEyCU7v7QLvXjXvoXTTq1zZL/EyU4Q//hPqkio
kusoLfOGSN67xQBBlVGY00QBoCn4Mxw2XVoz/jQACPvaK8DSoDCRgKilc5fK6jf4PXvrSL9cc1NN
aEBm3FCmw3BdYJ8L1cwRx8qDMD//wBlg+wbTzM9aQfAYKq1CeNru01iK7PjRvktDYq6bIL8XJiM+
yBu/jR8iaAQARMwO9dkz0atmWqGvtI0o2iV5wmc1s8zqyRkmw9XJ8iEoM+/ekTIHS0POmMPlDAX1
CSXZeNNuIJOe9emLptWUSzGKDYzK8kY5mcmjjFj+ur9LYo9fqkqIYeeVVAHMxtLwFii/Qi6S+paO
gt45N28xjRcFJ3eKzTiGYrZoey8vh9Mq4JrT4rvtfv1FqdgZqPDVNF7R0tK+u1hn6Zcye3MrPYLm
7JNATb+BtZz0UAidecEDoQL/hrSsR3vdKPbK0ZxKQsntKJOJMtbv159tr48uISfjw2X1RGuQKpd8
oZob4Yg4n+hKxyXDnU+bClqv6ymEHicyXIbPqs0GCRENbPdG2Vds5sXU0VNc9eh9mS0/wrCUmsNk
S7DaX63TTGA2U3cUVo0Q7Cm9a+6rseL4DqkpZKpTQthEbwsCZ2DGYpJ6eq9e79RzfSMSdLIwXCzG
5/VXPKXSqFQdf7pOrtVKpRrfoTcJLjOGQVngNYHByo099yXhF7lfrzEluTta8zeA9btnZkOdIf4w
I49eazbvZFw35TNkFGim+RLJHtzaaqXZXgJv2XBv2Fq54rzuuTt9k6eDxjsqcb7UyjhBnMzUYyad
gINskE+IEiwtx8X0fj+JOG5oBZbe+X7US8g0L52O12sbDBjy8GYduewtW8Y3wkjymOlMDvI4XucS
GWL9Eu1i9MUpAWlCu7PCd7uVha7BP2Ppx89gORnhAXnmA9cYSZfNbLLiGV6aKL8enC2cCqHzaaBO
mgqMUpV4VDlpv5PNoA7+pf3N0xqiHkP0xpDBVmh+mUiTRNE1YKjpTRqsFXZKr6pPRfxXIk4hAbCy
IqsO0bNetwFtIZVRIIow3vMSFZ/T7dAvmhlDd38tf0Zzkwnu7GOlEIr/lU33eUaFtKpBdhazBqfc
9YdPvofUYYiI4B3llr60cXBKb3rvlPbrZFsWsVgseTgIfJuQ053FNHQslc4One1bLRdIKIclCCWh
SByQIzulV7IvLEBqD8hl4ub9VeWvwGqa1aN3HUA38ngi+xA02b574YfE48NnKwfo+Ck+h2jyHUKR
YHpyxDL3Zlfbq8gzt+gp1alak3RZpLxrbV96oPFVpy0zeY7b2L878WLdPk6Z+UExszWE+6m6GOmx
KtK6Qrzjlx0pFPU0THtxHbswBhR5Q0v2BYZiXWxX7RWLY6ZRmgNvsxa9RYROvIZZd3B0hYIvNCiH
FNd9IdDlepkEBfCZuDmVD4uqncr2jGBtViEyO2zRBdafzAtEbGRhfztRdeTSEoqZ4mtuEYWSYfRQ
JkfmXI5qu+5B5+JXUWBluCGpJMtTGSV4mugMhiptDxnUKEM36OkZbxCpR+iSn8fVjd+IElqlNurF
C433BTXDNFgWfU4HBS5UxJ8wUpUUMmn8ZSsR1zw8G8kVdka6MYYkjHWiV2wNfzCicbGkl7lyOjw8
xHsOTmKSZYAmsI7sUnQ97nonr7UZ7IfLkwDcmWO27zNj94epHPoKVxWlei/0wBV5x3K0H3xVb5nL
whvkBXNZMXBltxtwE+QeoG3K4n7VdOKTxZaFOzGZQFdri3084VMlgIm4rCzZUFZIDDFlJB9BaEm7
37RUJ50Y7OaTTYmQjGW/4UDg36yhCgoIjJjRufbqXAckCDui+6vocuO/4suFofk1dbPCfwUE3ZSg
UwNqzlimdphe+fdFtnIpUH+PdIoARMwX5O7RMVMFSPZivdJxdGgApEfjvx8HuTbMrnBMVFMD+fP8
gEGOVBe+UPjo1uxgeiGvxdZzitUtRuAsP8ospg5w4vniqZwnbF8PY4XRIAuMi8FtXoKBylvRsBnD
72RgVTdBhWuVvhTW8Ago2s69M9Bw8ZeqwTjho64v17WcVngXt9Pq0nIuhJdTNrbB53tw9dO725nt
+iSMqyidxbmflrRHTQAxfvGvrbILycnc/pfFbFGfFnsI2Hbpmsx5BCluzyt4W2adJuMXhnygM7y4
9HV802BhcFF7IDFwy81zSi/vRbIv8t/LZpbk/WIo36pp9p1S+qsekgd5Xb12k0H0HuPKwRdA5J38
wW5MJm5RKEMM4jfEq/Amzi86iRkaglaeUcysUnn4A1m5MRxYU0O8Qeym2kGHjeZh8myRHvUV4/Bx
kAmos6+wKw2wcR0Id9O1HqhG5bbBvJVIVld80mexrzRf0JuORIl15PxrBmRKWEGQgi5jUDiEita5
85PIfPpRtHbNKDEIGc4gk/UE78PUxX87eC8LL0lJz7XY6S/XObZZsuEvNj7jObCevBksjdXnKFW+
SCFyW0ZeK/5U6RNaomubo1k/8yqzr5lfS0c3zVdXkzeI2oHJAt62P+4EsYblwPQyZxx08juUobzj
QxsPebfc8qXU4IttBrOPixiFaY+3h7YugP1uAeJbtl93BbTojNMbYw0efopiqVz0ZmIN7QGir9sS
KTTNKmqX0iL91IzS3/eJAX8jsI9k9sQ3q4kRVIK4GiGP5ny46qc1/fcaBEyG68yjrbfxLldV92uJ
UiystFBcZhj4/wgeOOm3VkL1nIuiIHOwJ3AIZORcTVyUuFzBDntPnBecPQqKk2Ea+4N48KH0MOH8
OH52wvH4fTx7OiQ7XIVDCLtpyV9Uaj9of/Zjm9WDDqVVuVIoOQ9UTda47QviywBx51rqn3oTRmeE
wj+Y0wK1YrjFMX5HSvsbx+jGJ6KgibI4aflX9piDS0dEbUJDnv1RyhJubyM1FNxmfni7qfBLCyhM
xBdu2qsgFKFb1cuit6AJqIa22B3UeigQ0C6s8aI4aNonR48bZIOcecxAWiqvX/R3t+WP4s03cG+Y
zUcuLA1ZVauSBYvM2xugGbnA0MCUSSq8I3hvmV1ikN7IhC79hghGab0iXhcagILQUsrzLzjf+DmF
I1tRIHRVgj8Y44eN4CS8s3wtE0QnKRq4+CaMttrSqHrery/HxGPCIvSH1pRA3eI5rAgubHTKgpQO
1i32A9zguPbVYrPQUte26pWwEd5Zkq/M/mp4Oohi09AWtqeeqqhEu5ilv2vKJZzvphxIjbYDhxu2
D7hWE7OP/AG8ZSbfzBpzI6auG7R2NbOoZWSCAB2ldyKmwgqw92LLbS0wbk9QJzgAK2O1qzTJhTVj
DsVAGphtz2+unyZ+05YHxRcP599WHtlJ+sMv/JIy7QBeRIwywl9zHDx8AgJLdMNYBn8PVW4K2KGY
qPlu2PEWnMjAexJGsv8+ZIOo3mOnKRAeKXXv4Q62HeiEVH21Og9UYtqeSqlYKJcclDdd3eJMvrrb
r5lRuq22ttkd0BgstKktH5/u+D+DfkbMGWgHoZgR4zfzYNHyc487OHzY4dI23Fcglnp0YTTeJaFn
okuGMxEjg6gLpsIfsTpiy+NCS5hlt5iUss5YIT9xo8J9CRnv0gseBVOPuCKcjRj9ji2OnKq1uB2E
wRwUyQYuUSW3TLEXvRw7rUTuC9FehrL+JNW+K6hMDQs5Czz+fUnuQC0GZEcAw7PjhT8qAAOOM68Q
tQs0zEY7M7tpb8R4qBQC2Ol4w8epCQApz1U2vIxjNPNk1J48hymQM1KTofzqCJSbzN5qphHkj0n+
Wa/bHzMRCM81NArEiqVY12WCVBJShZS7GynNf0RvPAOYs8Z21n6G/DJ8QYsxgrZyNwxezUZAyEyA
7esipEXVjf6HNJidO1sbzTl6OkgGPGoy9d4LGh0vp/2+UbSuNg9hw5EvJa8h/a/Irj+jr/ACcqu9
bV+CIfVtE/G8yS3sFSHL3zasYLyCiDXVA/thIeWn6TfyzvJhmOAXz1BgMfE2sj7UB/rEFc0scH20
RT5ZQ5phv/RC3TaPbzVjwnBqUtB0XDeC+C4H6Xz9wIDzVl93ajDrceWtXjDp7bjrhZSI2uwCwDkq
sL2/PiTll0Gjo1ce244DoP17ZFU/tboO4IhXPQafFsE3qKmFZ7X037NxPqkANzT3giU3ZK1Xqa4x
ziFB/g+55W0irnhxUtVu7GdZjK4UXbOQ/69nfjR+IuPrIAbPbiJR1hnS3G0jFXZJ1kK4mrcCgtrv
WYbWdy2aCBeaEvEYNWInLk6+IN5pw6GG178xJKypGgoY+eabaX83zB1jfO/6scCk1fc7DZMsx3KY
IvzbWNhtDJDkAWxHIckHuwKi6Ri2TQmu3n+zPFHTakqT156aFV48F8fAmv45Z8IM1ZfOs1R/IGHg
Ctl3OZqyhFZsTo2VzDrn3lTT8DPRWA64jwVS201TiNEa6v6mHvPXZrEFHTXu/gQm9AprcOs8F57v
EaMvtKPm9dnAOfE3TbtOimCUqPgHOAD5O409+1z0TxP40NtgaiBDiNjh29PqkDtPN/nwaIs6KV2R
IwlKuqWCfp5uvIrD6GzpbQsWxLxBYT8AC3rWrf036TP94Rv81naeRwUgH4VG/xrYzYCG5PabJi+Q
LfB2lDpUDSrrap4tHr6lkiwjQziN5THph5XM/VSNyrZR2AgqiapWgPudtgXhOHY2cQJVnvdpGypM
8UZ1kzPTyfrvs6rzabZqgoo1srQygwE7mCWR3ikQHTxKGfrNMIdg9Y8LpmNpQ1qX+8HZ6PLcbJFT
wsyFHmxLBiaqKYSQiaqYzol3K0r5xll7SQeTUJSg0Fg0gp34FBg/h35MQf17No3Hr+Y4H+VZkv94
CvFtxu6qbukuIlaANkyb9vIDhZ8uore1wPBsxyYOkbcVdDVxwmBp6MKLXkCl/dgmtLtAgrtNOWjU
2eKe7GUVkzPQNDvi6OXPdxfH12/wM1ogFY8ZZzGPI6yokW+3fbFK2vkkY21pNPHX9GJDI8S6mag9
kD+UexKWNRsLMg0YB24dXQsqiTipZAI17rTYhB9QfSJLOsx7qfyfCptI6LAinDppxvd/aP08UmuT
K2p3lyvz7vZywOgY9gGSUunADalQimiVmuDX8M8N6+q2zuy64I+BtuAIiNk5bLLPgM0qoOR0kYey
tcA15eP8oEQJjQRZ0DyEMirL6s5mZzG4/pDMVLmsXUoDaYNKY2fSIyDuQCX1KaXtfXVH6L8bpIX0
X+jzty/Yto8c8rra+2OWFdUJZYdYAO6GpAEccRLORgT9Jk4e9huF9Hcb40AAyjLJHsoHCoRv71Fe
IC5ASlh/6ydJ0LWTgFrRz+idGi75ZLB/f0RTsjxXWn4lAcpUpFHPsNY1pCywLSZg1y6nTsQL3+yB
VnTNkNdxIHdz6CPzsNowopDuAKxU9Bm33pJx0fm8u0cwDpxg6Jh0ZKqR/+tbhIF1XQ76FWudjXjW
aJT8E6TuF3hWW5gYCxxN2B6S8ynmkc8GdfJJBozdjdu0jyld7nplCClJQ880m6OqJePL73cQkATH
kBL5SELs4jYvVqaSundoeeWQw5OAwyElA+uxnbuZUVLdeE+gNXgfxnWtHW8UuiWLuZYs0Exg2l3h
8oNt5rNjetBcTHkcHtMb0sycLfJz/BqyersROAdakm/rcewj/lvPbaz+XZCbip5zzJHZ284IMOoZ
vigl68Iw8I9Q10A2u7GDC/qJlutuMW6tUMQgxgoYushESBNzDp2KTbEsWIK/AGV7zF678E8fj6Fp
73r2Wuf9l7Q8/RmqFJ3UWItImiLhQ/1wBjjU5FZX3fGbONcAoT+C79ZvXczwovSjyXsfFR3AxTP9
iS56dCxNZF9gvOr776m/FQDV7fC8JjrgSfH4Z6J68OXztbdeIRuaCTg35tPVKc/0fJ2s8abKJ1XD
3qOPR1a59zjm0VplSx0OBvU2EbiSyRQzPJISPRa/CZGM7B+iIHWBEN7nY8aKM7PrAZEvnty7llou
J8i01GcW6yRcpCHPj0H98B7zahvnwUgDkx35W2X/3Mw0W/eJ2Dwlx/+452RRXNJeM6ybHiJidEJz
hC56s9ua6FWtNvsr2K3wZt4M103MFWEh8hx76KWEaUOyFpuZsQG4lHlj1yMqYIENeXpdKy98QnI/
VuL+/voGAS3IB/5TFHde801OGYWbFbutqFGL1vuro76N/AKi8Gu+ftUZ+6DejHhgTjq+4AwTicR6
ICMVZ/3ZdqhbHsyKW0mZ2MlXOr8LVq4v9IXDSnWop4L+7NT4qoOOexWbiIaelaakgnpfH758MngX
tAzbzUTNwUuppNePhFRB+TEaLypPqDJ/CG77JBan61DPBg8TYJwQX8lHHF+WNXxSUZFYZzN9je31
aLWeD+HhVFj6QVq1osyyVofggwQdrQXuwYsaPi7U5pBXMRpRhNugbQtTBfwfLSNrHhxYPTeiI/Ns
A/wQlto2l1+zcl4lORd6gQEIsSjDa3VykALnfbuDhdvEheYQ6zeGtUJIJracWnIx8siZwW9Nu8tb
YyZWo+bsv/FjripIunBhZWHc5JFPSAJn92418cKANy8+Mp+wcXYJZGRtPw+5N7qTSlq8vINrgWhF
iFLMKzQ6L2CuvADlN0ynv5nHVK1iIlFo1H1SokCpdVdVXGIPT/lmzBZOzmbbN7voyikylYg/VxGu
nFPjU9KRbraBaO8u1IVbo/60fnk6hkhS+X1ISl8h6jORn/QKe/JaG6xo+zf3lJIusPXLYTUzP8tg
ZVIIh+kxf0WjZdRNU457kWPc+OD3/LKaLkEO5Y8A8h6UpSsRwVNb1+p2+UF4PrxPm4IMrA6UE80z
QYcOu+rS/Cm8rR2Vb1yDQGTDlHj40X/YsqEHNWnLzxJYmn77CdLE17vi8A8/enKlKPVxVNlJlFqn
UXR5H2rPCAW2+nTozza62AxzNxyWw1X3z25ARz6sQthF2wtjH4KxYXyuqRTjJiWL8FSe5YwnWGFp
vJbjEqaxJolWROPy/CYr1fNmmB3fwWBzNoJUFxuep/5ij+wF7ejK06Ntk6CWh98L5AhTXph3dcOy
m7Zzk1tDRCIsam3UWhKdCqdUtsRZrrBIkAFTPohFTkFuapxmXptrziMXeeG6whnfbskF2JcXBzwp
HcsKsb3ZYmG84odyvchGc/uKCLbbsXZIIAC8E4MVMiXzbZWbNUpBWSeN0UNdqvtaSlUuHPjasoYC
norI52xka13I+bOn4/4fWur6vy+McKj3pWo6c0Ax2EKkd6H7tdJLmYabaRIsSRzewqYeV4icfhlK
U2x93fcyFZnISJYcWXJhir0HdhG95xVElantAaXV7D9SGIczN+6x5tn0NH6Lbtn1+1p/1eFnVU5K
pfsMJLcq446yA11FEuFE3dJTl3ZZ3Nj8M/02QVEOCGeZBLgquKqZb7RDiGje+oEBiD/PQkcUGind
DNE22gAMSwz+VjCQmBLnqJMkb7fTBOkfGhrLo+4y0/0rXisPFVnStdibZlAUKTqgr1DXObAhRTPk
LI3wS6nFsHgNohGFZ480L/ebr95si09FTgIP3Z5KdQZn1EfPSfyhPHPJ90vyZiO+xjtBvNNxJAvf
TwyLyldOTfm6y63zJLMk8nao6Iw0CKO0Cs2OuCdd4BDRqIoyKgxNtpLHaCosCTblP4FRxLVaYNTf
pXDqz/cKcQrFBEDY3+XtkJGoX8ch69elQVWU+NW0JJmfnDXYuqPkZ4ajgvgulXCxEY/HG3oaYVbM
0CYDsX2ogrpjmcRVSrtHLmuZL1WFh0xSwiwQ46lYXuZYTeYPvptO14FX0hQ6A+unbMpza8ss3IWz
ZaundAdoRg8I+sEClNRoP1SsdAfYQ23zIAANnf/REfh8+W9HhJkobVlMuxRr7BNVNVjp0MFCJryw
1pg6YKJNsJ8ClnhE8kBF3o/kr/Qs5uXkgoqH+SOWAv+XKtA96uKp2X3VxPhhj2N7ZYWtcdIL7lml
Kh2IM3k4YmhDVsljrLSO471xCl1UeU4f1GfUCApwLoecVZS1VFGTF2uXVDBX1WeSoUZ9lfhnGIrn
Isk+BIXo+FkmFk0wCDpcjUUeW2XUiXhokAd5rQCBV31KwlhRzzD5Rsc2UumGoIlr+Ysup2+m3PEi
beXOhvIHr1HA+sWIclSFUN3fnFDaVz7OzgfbpdFjTVdQpBgg0x8abiOLBHS27YDJOtSmesTdojZY
Ov0OftNVF9qLadS9Jstd2Ry4suj6TkcTIBYLyHAwh29xEl6QjSr2nvrLhlrCwxHRB23DD/0yQj6V
oECyjMg7oYNLz3A3oRhb+uCoEfFESVWZTeuSumXZatt7GQIEwvMLN+E3S1zACKVo+SGD/siQywyS
2kJGKqPRDuEONeu4uEQVcdbafA7rF7Vjqxv5Mh6O6JvsRW/UvEY7fXe6WSMirOHwL0PulMZqy9OK
ufTi+NaZN6s1HYNIPxmUKIh5FgAZt6plol5XY+eH998SK/9UKe03r6M9XLSDFpNjXSGbc4YHVE2N
bzycll3qIf3bx2vRPekowQIgK3Faj3uqK/Ide3mVuRoSMCENAIT3d3pxV/2Hdb7GFv+nFTTn+zOW
MwPEacKO2QaVRrPrm+gnEDVgIuUA6I+G1v9OKUl1O/sK+mUNBXVwiFz4ehZYDrJ/g4ntSL8Iyvg/
o6/uQaTxv1gBlIO1GLRO0f/bJ2D/8xhqw968Bo0CN/cD/93gjCaM2vNQjYZK+SMRhi99hjJo586l
3duICCDXXEmF5dnWtaZMBr2s98SmWRzJKdXmpf837PrAw8HuCOeYnJN8jZagCrNNaso6W1FKlTRn
AqYZfH4K4wnVtnCpd1X1/oWNMOH+sU8IoUlf9AuWUfft9xC5YAwfJHtu7YMua5H+noG+WCUhqhHK
oQ44sUmwrtgmm/MAkSCOQtwZ9r/hHbAy8ni/LeIvKjCs1U+tKGMXx/d962sT3vh2Xb1mZ9/R1QBv
JYureKr/GMOKg6QSyui1Jjm7+kVCJ+2qBRDEoi7iZW4uUiaBKo16/L+lwORIY9pBN8a+YK0Yqin4
bNcJhFY7mbk4C+WhEABmY7KSCzR/rVygSSjS7GR6iKniArfpnZB+rdT/NNdMHppjbn+Y0QmAPDoO
/41Nf3BqNykQfMqoBYDXb6KsSKZAHo+icR5ubTxwAGIJ9/b36SgwDzRfYtBGhiN2ADvECawZpq1C
aWH/hGJSfm1Ah5cfahAOetBF6vtgXFkcxHc7wMfxitN2G1oGyqYXPdSyn5tr9sm4GsWT3SjBvcwG
hpKXtTheLdX8Gfhv332LNC7wF9gnCEwPN4S9CJCETZr9tME/mrFtZVqrf6jYgImYwftsVeKqnit9
vr4St6JnIH5Z5vIuA7e4NMvgtI1afnFB9FmoBqzfkoOLRDBiVe6J7kPvE1YDhh76Xjy6vKJOi/bF
wKu/Z8pXNuU8Qa5lSWjr/X4PptgyeZp0zgFB3F3Vpj4XuQtoskqCd5hLpgP9MY1snHgTkOR1Iv8d
2jwzN9hdVfd0RARepueW9NbSUPi1t2sN81JKbU9PZhBJ8r+Z7R1hVnpIfRuceCcfh3ENJxef2qfl
9v8GjAvnI3cCIaROWGXfUK/GSRNWdU2naNNFlcIrHFzyFO/EMkC7pTMXe8GMwq08HRoTBsanzFRp
JDh8iPjViCoy25J3JLSThJou0OUxI8sJARXGznVlFDMq/qKdTjpfV0+YIE4OKdzSNvq48nTgunl4
v+x0oSnCNCTtZ23RIyIECaZE3sxN2sLjOf540ueWA0Xs+T1N0ILz0x22X2XaZjEmbqRO7j/cnCEx
kr+yP/ADP186+BpOFyTDMnJ4wTI/J0OqK/h9+N+HNAUBBK6FEqJ83bIbFsNRHIItRU6Pg9QbVcGG
zrASJVcGFS/K4vfYmImJQR4KkUZMGQzxkV4JirfvqId2tylYcJTNltu8VCVHNpunKTATwe6fdxje
mhday4pKw7UciU484rN0sxo9AtfvWyKwb4l1GVIBEWGBemdUxOgYlxbOppOA4XrEz5rxQfn2hBYo
yJRw3MjILQAdI+FM3+RzN0ka4ZxVPlPqRjt2TxtAMiGau4XQPpb/VpTS20GGYn7AvUKOb6FolBYV
lWUmj+tYU9huhjZIkvyT5QSVm4IxGvn52isEH6/kpWthdtxkvm0vrN9hulyMJ+A4zBBcPsTqwFez
C2KY4B4/hGztBBiApbB5e0hjiCINK5zp9lkYly6xR7VajZSOZvLJ39BA40dVn76Xsl3ga2Fw3AOd
tWOUF4jIOI+GjGMlFElXXkleo8t0UwPY1S0Xe42EFg1YdmUL97XQx1AU+zxrPQ68VBcQXRjh6Tno
CXU7706Xk/+5r6bSg/otdza8H11JjosBJQjw497u1fC9n/FODC/KmIIAUxnwNErBMHRin1TLvxfT
PCxwafrvXxxDVap1tO4syt2KRJha7XodJYLi5AxN7CFayHZ45a5liwHvQ816B0U7Ej/KWprJk2s/
cBCDmi6Hc0iExgW8ynr9PPE2dY6FCsCNMUZfofaN3lK9p6mLbSmb+tjgQgsmnw24RalTpBAi4IPq
TsKO3S2G7N6npvnCt+TkjnWf86pek5oyxbwCqbR0IqCKXzCtvU5UqZOWWSL7JDbyAhrbmmhrdAGA
1ufFnw3F/1kBbdpzwrVcZAVfzYrS0o6AZ/D2aMpj/kIF039CHd+FKVcEct3ylF4pKHQNALKqAR/j
zd9p/DSHpOE6Fy5OGJfUeQA5XuHdMJJsPbfITT/f8Acxu5Ttf8SWfI53HhNffI97y4q7h33uJplv
PboEVw7x9njJqF1Im+U/RU8aXEzXWODmQtSXWI9vF0wTOBgcK3TM/KjgqHpaU5zyHFov1RnoGcC+
falzc0JgXTeUwFqXHet2I60eTuGtV68gk7IgSoB2abF8rDSz0q8LfcjUAuSjhjj5jyhDkuoTg0p8
lWA0Q7j1NtVo7hIIBB1+MYXjYifYMSdbQDgfwvVtLsEkbbIsYi13y8TQJAo3ojyYhYfNnSQgkhkf
Bm9Dd8Ff8EhVNpL1J/HPc2eosazVfImwqn9NL1iMLWtHLp2qhC6GB97FmjJp9uDUeMc2NurgMq6s
82YzPltyTeoi2rATWbdT/frqlROCUTiCEvSq3DkBqeHIabbbyO8cXuJ8UdVHXGq30TwGm1oxXOWL
iE3Uh75J4qDLYcULngBOlsApwJ5d5YOS8n34v8yycRS+i2lOgCcrB+wNMwtOvkE3kTm4FAuH2W1U
H2/PP/voJiCWzD54rPkbw0FDBk6JuNw5pmvMPYFgNkcu4mQKh/kI6YQQTh7G+aJ4yugDmilq0u/y
GWp02J2duqzqdXRgHG6fQ/EGkUaVufSjfDpAzOy1sr5XKmFabNdLXHlfG4arm+pKjSqGsUz0iubO
7OjT+nTDJ5JoP/W0PSjasxHnFw9VRPNqf5gXwvIVr96e8beGuyC4AM6Acuen2/EzRvxmZ4k9SvQr
xHijXIR+YnVNwtEGg6hnUPSKcQNjeLWdniPtBMvB7q7p6W474jwaEzXXfp7L/UxdGNpllUykldl2
GJfF+e28Nwc51kcNN9nbZTtzZb+T2UY+3dHWwOLPY6KJFiX89y85F9wPrst6Z+f+JAyKR4BPf5hY
p/wffS2e0rA9FaszeOEKYpgah2INj9AGREJaUXIVM6KIsSEWJd8ASPqjO1ON8FiR1DSXiwcCRfte
OIf7nKR0T0n6wdWUFuQb3zMPsp9sJFvFMvMktSi1GycqHfjyohct2Bvh2bU2JimjXPsMizlVaXjG
JsVLZ+GAesoSgIHMAzu+aEIRkFfkQ8PT81IWFcPp7vH8pmm/XsXXXXU1jZ6XthxBs0qkOGJilrb0
Egrw0an3kzWY+2Kqndymm9GUJD4fx+oVMGROlRWc3RgRR+dTNuk+gzElRE4Y2V4+PU+7qVQqHtKn
DZOrBLaF3btDM8tsRVdde2CJkeF97wYJHPTB+MrOZnIFHIn1IUqA1LXNBYGTaf6yhdzkBQAgsMWv
KNOvSGVIW2kQ8FuuQG06NYRmfDvWQSsvHB5oQpw3E/nksxMoy4XrgVlqh6htyqe1h/096o/EGrHk
BadoN0DSWQhKwKUKulcwpWJfESqcUYgQuUncqFMnaWNTC1VOt5sELTMztxMIG0a71UsT+dDdXGEa
ZxvAY6m8Awvji4nSRtIr4MV3l6BoEmNQU4cdVaR+MBPfVVB2afItDPWv8/dZHFHwfRMo0q8ryYpv
IyiK/9DjEZKo0vLeD3P+FHMmI+vOccEdU/bnXbgyurvCDX7wwX0o/3PUE4jADgseAXXlN7yt+Api
ezdklcQ4AgkbCf0teUyEgOKgw4nGLtRt1i9W1KeMxkHllMnoS3wK+7ZKUP72u7tOlWaOTmMsQyQ6
bfvpyYdHRwIbgpOfkLorP3OE5KnuwUTVgJaig0AImBH5GWgbTSN5OJh0RxOzMwYhufMGC6EP/aI8
7TkojeiDvJwLKNywRKcxNg3UxL6/M39+FPDwSYSBxD/7zYbt9kM6r/LqaPO3oRUc3/UyoWXm5RrJ
y2eazIO1aBLdA+Qa6mNjkGq3vb+a67kXmjI8J7bfnZwdSWJ8/cptCVIzRp2sDFRFIJJ4i5VxGBWp
EIdiqde97k1ofXfU9CYBYNvrtAxL4w4EFuP65yfqSKSn8cuhG2A4S+P8dXMH147NVfQq8kARFFJZ
9gjCYbCn6Hz/cxyqkI2VO2ZYr0CTdKm9MOLGITOMcYXrdCA9SYj6zoP48csyQE3BHqz5GrZrWiif
dI6gGE2xfLH0iP/y/nBD+uZsfBr7q5m9pe7vdbvm6FxWmN0ElmgAhV70aoF4jIGRazApaWPvGoeO
rJxy7yDgKx3tEQjc8kEO4uq+q5vaMNfA6bzagQ5Li52IMIKcyHvun4sWQ+26zu5sl8Gpao8vFjm0
/07mvMO/yauMRiU95DRWtpYxxundNQl7fRcpsLa2uPAqwGJjE07eta+v958BZ/KyMdXg/RiZYuoc
umY6stoLtXgDDWqA20ui52W+Qsbj+QA4HLcGZ/F0LVz98OmO35s4uhbpgGLosir7MiH6glYhYtLi
B6V1993weKCKeOyGYGqFbMDfi50Bvlyg+q363iDLYCfA2RsgzCrzyOt5N/e2pBgIIN8LatMAkLUs
LMvijFtggSjabezDozxlCRBdZJDn8EA6rYOop0TjSlgFm+GEO6Te4d74X0tRamP4KeBUC5FGsqkH
IkAL9T2GeDXzLJv2XVdQo6mgqXacbFozr/nytvXyBlKCYC+Y66LVsXBR7hcG8MosED6cG2ssFzUZ
MUFlQGsKk9lepAMsk2jsT87uOKw0LrT3ZDuGL/XYFdj8NZJ1vm2DoVPzfX1g7A1LaNEIFCyq/JcN
Xm6feS3NUuwq9pxxhYnTs0fOo6hc7pmPkwLAKHSr2KUVeMBMw7K/9qb+pOSRfKZiJBM8y9E5GoPl
NBbAgdYSbBYxd2BS6YOF3tGkeG0O1dy5hq8Sp+R15MKELzactnODqetP7bNUx2mrO7+afcKW6+Ye
SixqUWqO4SW+NlQ8YUXL2AiW4IDGMlXHlqmmzBXMoF9o+0CxbeBDoP7/U3cVuPH5ks5DLRdybbHQ
jTgcblfQlI6R7Y0C66Z2WtWS7SWDfXrJIU+8J2th2IxmgmtgupNY0HsCFYp6bC5/UA1ZvXTsnn8/
hiBM9VtTa2MkhleAW5g5GOGRWMRQsHIAF/L61eu6iA02D2ru/wBhBlQLleEkzz+D85RRJRi3/f10
afNRh9dfhn935YFby6QytYU9rfJbn/ybJcVKVG754zka1eMW0duivKszaFVQc2W9AOMJsN6zFHBH
DOtplz/m41SvyHzWHD9lGChGz47++v6ZGvMNU2xzFjtmwUetBnQnlknfKaulfOuY3OUjVvoXQ/jU
SoRHdPyFxzCaZyGI/cn2L5wZVbwwBFh6yZTaAzVxiOoF5odFO1wXPmf+cXVravSJPICRT1F/pSsp
OY5oMOtztPJsz7EvrzRBnhlTNyUFmpQD0RSkLOBqZnR9bORYnWtNNKNLwHYCb9KrJnslmIhWHCRx
9+JbIsVPzAfTZgSegI8jCnAb6MdWxHujNiFcdywcChWPRYqJbLfCf2/GdB4KBoi0LXTraTe7FgEZ
ZUiJLtrWkG3MTsl3LzL/9ya5dSMw0CmXcerPAZr5yNJftVWlqXEvPsdZmwwKFCTBizY5ZJvmZYCR
bahEZMQzgH1Msj0qxxhQ1XKzLZFUvB5/AFRM20ONnW4Oo+g/nCNV6cyKVoIWmhfVZodju1SE4qAm
sHyg726bokzcK6ooEJaPEJzxcfkevzw0iHykE37UWfn/nlCfGzc75Ih6RqI8Sov6qc0LCabkMelJ
3NsUjJFKeKUv7yGLPwAsIoAEi+aOE+T7UF32Y7w6+TUcEQvjMIQ/Rfy273FGwtu3hkZ4CTgZKVoK
wjGGEPhhxYF+bGeqAcEskRMjcZ5L47D/6Ll3PB8d6lA/e1uEwMdHEsR1gtYcrNJ9a5LNb29zQYSN
2dc7USLxfYgbTU+mgxYQ5icSz1z+KyNWdrkrrQ6ZwB8ekB38hZK/zWlb6p4i8yM6W9dpzxk1rcuP
W+wRMnr+6vH3Z62pZHAIUPNGs/POdTPRzCmOjN8hu7AsC1hkH3gTbwRLjdQKM3+QTLJq3TE89JYG
UDuW2NMbDB6HYiankxCm8kdQOtkabQWHdlNtOvMjUXLzX5047WRDRViptdwP+cMX2+xwrihZpBNp
o/wCTw4pFmtiHrCyQpUhNZWEgQXROn2utWQkezhpA17AGI2zqZc/Vmee2kN7GuzqWaY/fMADnl+n
zpv7WSMKsO3MZ4HICpZCQ2Iecxvtv1VWgUmdFXFXYdIFWP+5S9jQNYB7K/pilIgMNMLZx2fJYTd4
Erp/QqSQQ2EOyCxTrjAoUxOHx1jpyRfcSmkdvKB6G6ZVeFdk1wS1TRRyq2ZyugmoiS8HVR5U6E6Q
JOUipuhoxiEbuZGIw2pl6gSqwd4It2Jz83vKCqWupHqKPSlbokvVeOcxMnJgG9BsTUWvNJko1XNh
53BNZg9J/Ymhga9bwGqM93VqAmhKFymgszCFTY9XcQ/TAWTocDmBYbrfvyncq6nKzem94uaNogIn
uCGKpVBj1U4nroC6O9ljL0i3gazY9JsPIOYygw2r3IZvnFhTb5prrnWqss07noioRrgfCtfYPxN0
TADRTd0azgVHAw6t4mO1SW2Dw3kaP9D2A/tw3N5keqxnjN+2NMz78d9NUQRxnkeJkHtPAww0U4zd
SxksLH1PNypCTRTW8MaSRi6HbfmFaXN7O3g6UDsvzKngxyCfpzMqYXFizUu5iiSkJlkO5rxNWTYQ
BmB7tY38wedyMKO07ZzBYR1TvMUCuFGCKo5R3e/tcrub7b3i4JpGYHF1OYmDyrMgwiQLpCBu2/NT
nM5s/IaL9V0MbZz6W8DA9fgdNAvqv/0oOZfin7/+RDqZ1G/uyqxPHOlhsHCQO6HnxKqYgRbrqCun
eV+xMwRlwANlEZkCVq6fQUjVa88asMIa5/jZq4j7YG/dd2SHgbrprGAtZX1Ca+AitRiVyny75BsC
8XuKfnerzA5G3T/FpTu4gRasSdirXamqJqWucg6/caOAGy5QllinT6/nre0wxaYdewfxmaIjQiuN
VCdn68sxqjmG0Uzit31f3R29gqPVkljeEZIHEEbdRuEvrRYf6uQ8Y0KuTGli0nJcx1rLianpcjT+
+sNOlG+Vx7QrLDewOV9RIbBs2ku88lrg9OYrd65PMa0yJlGp1DDli2pGVpYoXXF8r+alpavInmPt
jBPI0OeMDgf5Lwh4vQIvOAC2jb/j+/7qwSq6Oc7/fybW62iPUOrak8ULGJLU0mlL/j8k7xRdi2l/
FpTzIwVkrDgGfxt/4CCdNRgI2vWJn/efCoFfEfCyXXPlVQhwJ+7eSiZP81J3dGKufZF/miKDGy7p
AsWBoixstKGCzgt6wD4O+ZamKDWtxy5tijn4gn8CM9uRk8wpCnPu2N0+FniMtJ+K96s8Dyq+Kya+
HLkKHKCP/90FSJ26FyhUzG/vaMYBWME3hLJNPfDTA0uwI8tebbuqaMXEf/591oh18yS2Umvlxgnv
zCdluxx1XtQAerJaOv6skUB6JXjC/WMta5UJOBRAmKdA5RvecN6qF6e05C1i5wqqkGhgc6ow0AMJ
tDK4PNJ6KbgYfih5lt8qvJwMHH/qXW3r5q+GLa69wp7Y5qGLRAX4TCRbSoI0G677q4+eKqMzkzlr
fzngVdomTtzudhxaMF64fgkP7MHoLI5Uzrn+muY2nrDVrjFFly/DU72CpBp4hdodDfxTrZQGob+s
cwqHHBEuCWy4NtlMtFzrXlV3esDjLhYL9+By5Bji+o23VfOe2UuEpwhjlEcz5jFQaYB+fBsbl8vH
GL7rXh/j1LaFaCJoDXGZdCIK/FwCMXnR7AeAUTst8iFrki3wVCRsVsxUuFW167oEc5gUJqWZ5aBW
kDKQpFJPa4RWVuCzOJvJiW1CHmBTLcMscF7wmzhefiCbuWifdnfPeM14uSf9E48KMfVJwgEwfWYc
bNeM0f7QgmXY0ydp7HYEJeDQTwr7ownX4KoOAUI4TQR32P7CIXOQjbN4nYZU6ICTfIe87VQIA2cj
TJVPN1hOlghKQ5Rx5MmleO2/wd0xEUgcoaLZ/SQGDxkVf92bjYbXHpm6LAcQp94iw8i0mtRdajma
76/rjSzHRF05nUtjrF2hX3FRPoVKpyaxaGFxEuVJM18qWHyu6/pI/BJYQYS1vrinuUXYeSpt/wTn
d/c0GOqUVqZy4Qxrt0tMbYazQWwyp76V/0yDFYTvoP20vjsCFCZK80bgjSXpj3WqWrJRxSYtP6lk
a5YR2m3kBJUqqN0t5efNULBqYxT9dNKRIds0dlpcAPHF0Notu5vN+P4UDA4kNhVdExRhZfov5qK+
K2FtWYLiFVmoNzwZ5YduQZ4wdB/E9sXBRlNn21IxFeiEQg/Gra2M29a4xr2W03nfpU6SmbgE/240
2hurLR8tYB1s1gt4VpZPfWKKdsVPkO6pY/N3UoPKJJJRjFLORsT3q8/t4iguYjE1kFb81VS+Xu7c
qSysFCuu5Ytz/zKSPSw+4HyJGd0iMt5fKL9mOT7BQqaTKjLlNCUjCINIH3RVhoalkbr6P79lgrwe
O+Hlz/bfgDPE5aU4DBmvnGqJUGkxQdOgmsQdN8pCbVfiOVCdxXXEEIrNryIbNEn71kQ91PkkFzW9
dxiXVcjATG0DNOQqia0Pp04H7F8VDXyskrq0fqf3a+TVGq2bIeU0inJ1fo2ZCzlD+fG7+uEMlVUQ
azRuUYGNynYzaScBiPP2uyTF3Fh9wUaTC3q5kY8HheElommkbIqTchZu7uce5XfLDLige97CuOvc
6GAulkJi3blMwJMSH3+WsDfSrJzB09kV9MoEzFkLrBtzuPCHC7Kfb3qdFMvOqGeSIcAFRpaleZ71
brji4mkWmbv3vvIGP+MWXotdsvuariBZuLEIDF7NyJdIkjNbLQGPp9fNNvJzE8UD6/bKCx4m1dJX
/Zt7OnC6HEnhHNcF8x+jcRT5dVTPNf+ebi1lgzbTaGTi+MHVXarZzdKPxtGvMuturG2+8K/H0InZ
/1x9+PK8ntpiJ1VYRRnNI5CFt7YDlY8SepjfzKZAxxe9C56nB8aCDoc8fKttxofx5xQqV4bAIeNg
WNNci9FHa6N7Lx8q+bgRb79qSADhf0n4bLTB6baJcu7YDUFztzJNC+sbKY2+vYa5mhc8u8vt0sUA
y83Nvud0cu9OZYnb3x2vR7iYnDHBRxFNjBugbCmbCBSTI2cyFUalUpK9nAqAFylvEC8Mn3xGZnvW
/VrYfh9I/d3E6O9UtsXgNa3Ts2wBvWUV1OPuOKe23cpyel87BKfA3YNwawV4wjv4eetaZi3/T7DQ
vrC/V9PRY4TtZZ8bTzjDs2xWC2LOq6MIPRdV6ua/ueZ09uEzrBetJm8twlkYNmbbOedjI+8PmSmM
pDpv+GaNf4qVfQWmM6eOMr3vF8yoUttwrYn5HaMbU1OxNY6mwhWigPgm0he+nfS7luxQeFtwuAlj
fXtGb6qYehxKXyWITRbcSBK+lmTp/9EWvZzfVjgQCQ6EfJ0jRKZYCEo3vDsxVOirhs25A6CIEiH5
A1YTKcItp3La7ywmydj5wKu2fQn08RGY0uX/ZjOCjtC9i/cQ+00LzaTIYyy2eoc15nFkmTMqSlxS
7XpqhurFbEa2nz8nc4CJSpnPRYn7bbMWnsp28HbM/3LqrzqvXCR6i9Tbzh+BuOD68C7cA4inbOSW
k4SLq83TlJkYrfSmCLmTKiQxMko5Fdd9ZyL66n+bvIYVwBQCSDuOjfWJnZba6jxDPTD/x9ExzyPc
QIRv+WJwQE6Rxqai2YKDV1xCBx4Oo4BQzjqzLTtZAb5VG5QKylpvsgVqL4CL94D5/KR7UIJ4KMxC
NyqpICJ+LpbXJg68TySVtoqKJAkcoKIelaKKWdexarjY3J6tWgD/lu0RngHvt9CbzSqui9SrmG7n
Z20omDacmFhja0WGWvkKSxhSZ93ojRSOU7Tpd7buyyd85RdLWgVQqU650yLtV5CW5WuvLnBls4r7
I3DvnI+bJEPt58hYBwensUpsHM8T7LV+HjEGw4VoSPy+xX7gKAUGv3zTe/SsoZ/+ZBKWJyVOU/ld
YcaLzteZUCKzMsxLrsnprE6LQQMVFAilnuaWXiQx83evf3tStGyZ3PZ49minW1hapESvqV58C2Qx
PcNFjL2pco5m/qK+Q1/W2kGKcScJyRwlpL95S34sqy58qhFd8UdNOp3qGOsKfZg3bX+83wlQS9hR
d4GwRJZHhUEG6WFHSRLOm3LjikToct3OCztRovqk7OmDSd8NcMaIHDlRUFibPrTXWDuLi98vaunr
iuCVnGN5ghSuwcCy9aOm3doGqmYHlJyM5lC/8fIWEXefcfvxyBDrKqxJmdKxiq/+QvGogWQi+zvh
Eev86prGGIkTaRgvcfXAF9cbLr1qwzGTLQ2WI8TyPxd8pK0f2fKLDgW4n87SCQETYG3R/3XaXP5d
aA9/2MSfeaM63i7VaIAhkbKMgybQH5GyzrNWupBmbuPX1oOJSs+jq54DTecazzvZTplBJhZ4/Yaf
l5MrgWkQAUXR80pD4j4bICF5fQELiFenYEMmjG8YRQChsDGSpRxrBz1rTSQpTmw44+J1KxE8dXML
WKNuS6FXf135oPQCoreHMLVEaPGAUf/2J6VGP9s8pDlr3NE09OIyL/5pINMqncHz+g/p4JUTeqvv
5GtShv8MUPb9A9+BD5ioFpVxTNHwZB1OZIqznjzmua7hWjHxVDZmjxB0eAKDbGyKt6rxk/S9VvTk
6D9Q1jmwyLtEMQIaLUu3SdqpB0eaqACxbAbUWAZK0mgEOuLzsNgjvm7ocF4jqlCddHHEs+t7TCuW
oLqLsv28DWvzoXEFn4U8TH5Eog6KpyN3GNAkBNH21UzAHe/v6F0ADsgAqnJuWP8Pe/KcVytmljDX
Vr4803J1lnCjpXeA4VO/GVjMaxgiqJ+ShazMUjfxBiGa4yt8rBM/ULaFz3GoW38YPDUjizEA3+I9
/Eiay2iOIYoPgUbPELYS1dZvkpoYOlDeXuP4KUUT7iWxqatH/u/4t1LcWCQGAcu7ROSh3UZfSNb2
eINMc+1vpQv2HuDQ0GOjtdv8NKeZ/U3RpgI3lYOvTmcjXZUDJLnI4rwhZYKZdU+wjEr3QqgvenHZ
lz6vtPkFOEhiEbjg1bNhqwEZWskYtfTmAvtN8a9D33UUH/51SPhZ+QkADcHWo+H/papuyGzdLipR
1ZCIzYOdJtcov7M2xzhwnveKg1a+yMqFMo9f35aSiUCCriPeZqUpXZizzY9sqzAjr1ny+fq5Q95y
dO3nZ0EHV3tqyVzL/RMb+bnI7on+Rj3WpUnmxr07F3RvMBitmL0YWXAtqZfipYcmSfpLQiT13Ild
Wa+o7MMOr9v9XIY4WpQ5f3hs3ugiv84/ZIiiVHB/JDZqhCYXe1B9wo9IDntvk90v4FQQsYRSCoCh
MwRbbjwpHBfa6d8z6iCSR6tAijbDMwTtNqjk4blSlXwWXTp2E0sHTVUeJlVJRqUguDFRM2hJejiA
6/kqcEq8V0hqqc3rAzsrGi1OjiUUYWvFI+dgGDXZ+MrXKrBwn6/kjFxsLutSviAzORH3iSFeHHAe
VdruyUK9+TpzWfnnj2vWK2GghXjJamMwceqOZWuHY2Jfvf0+I0GVBmJ9S0EPBmCEaiDdS/0sm4Ns
MF6/z4Y0wA2ggbzsNYUVy3Bjl+/g4XOnyeJhdQs8jOz5PCssjJFwISLGfJfAD7MxFE2w7dQog12Q
qn6I4T8mC+wpDFWOqqGzhI68I74XrDJt7Spu4D/ZuPiIMH/UcwBg60YPnb8EY59/Fjo/6TsX6aI/
ouG/Qv8hp0Yucffl3WIRUUuoWIp15pl6kVkUaCVXwd2nQ7HfZd//jdp53h1LNU7B5BuxZYVhDo+I
brBeRTu73ZKziC+CY8yhzExwrbB51iE0ZSGEmy6H/zdUbex/b5IsmIMbG6uV4Qyt3LzD+rgVJW2S
AE37WUXm123Ft+q9eknbU+4XXB4aT1l2104Jt9JBFaZLJgFE1NRYdXacTc2zJ9a6uMDdsXLsjmNp
h9rJ8yBPgGZ3od1G9uoRGvGm3GJnsWFWTCZfFbpZxuz3T6BxH/0oAYIyOXm5PmwotFQjQpOOsi2/
HXnGXVRIq2D/DQPlyoROCMhSwppZAs/fohYzAIKI9UQ/sN7iHxU7itTCxSV8BpEAf+CA2aWkaqE8
+rXqEWKGvWW4HkV/DFq1p2A7szq0CI2nlpc40oOnQCRC+Yf1HbnV4zylbr6fn5WrxK522Ov2egaA
R6UdR1cwgyJUSN/Fww1Llt6IIjPTfAqr7URGF4VN6k5tkHzMgmyJm4lFfgm+TS7aNEUMp27B0ulB
6gKph3QQV1kl8zedtNzzexyXypZK2Csmjg0xn52ojVWroShEDxDq6CQGplE+Yvf0N28sLmhA1lNV
4vOWiaL7CkpD2YaXgO8+5jE9mbKc3BgbqwdZYBAjShfaMNR/ke2MGXbth3LdeOaYH7a1IQVABOEF
I+YUioLXc+oBE1ZruArasUJO6100M+tiBP/RhjNX6WYzHpBSHdikZEfD7V2RQ255cF2c/8/i/KAk
pbDqGbfnnWuO8TULmq+REuft8prYPEDKkPeg1zuTN0CVBQjh+5+aNOTLdXJkBdgxHzybKgikceRy
5JiFfnwmX01Ig6J0S0oJjbnQITyGu2ISl9d8QMe76kc7inbn76pnh0I1erTmf40VNb0TUPU7Ws8I
TbHCrtNYsAiEMIQ9WR/wSC41mqKFqKZqZFcivlwLbJXboX6Ll25EQf2K+HQBGECo+buakbQcnW3+
qtw25Tli7WUsKaG/cqrQjHR8lluGOU7A90RbWA6ujB7ztqZynhVBEeAYgaIsLaVnMUCpY1KVWCgp
d2hT0d/mJBWvM8KpYgEatEU7NbZ6kA/8ENS3AL6M6SN6AgujpwJhuPuTqOVeIozLWvil28zzDan6
zmiPiBtQ2GoWCEGQTSPU44rGG45flzdy33ouinwxZ7dDy8ZGjCd95R0vtHxYIkiiSfsuaF5u/tDo
ebGi+8SewAKBy+U/qK4AmqaqOhd2bkTwLDlHiOFUjFa9Z9YgsaYXgmcR/Xn+M+Qd+pjy8y6Nv2XJ
6CZ6zITjwuS3zwGsQFS3TqOT1ZeNuqOlEgvY6zluUvq5GtkjudpQVkVi4ziuAGbu0vf7u0CZQTw7
xpPt96uG7MI1sf7dAGlSndp3e5GxZMNkxgC4AJ4nvaA2cvXJbY053zH6oKlIsJrAFStic24CdU+h
P3cY80c944JVqvZm2gg6ZXB51JU298jw/yON34DBKC+nOBgpfO6rRY4FPlNy/Hida0ssDjZH8pHS
ONkXD+gEfbNmL96zCXHvVyRoaLbKaElbEgUbdNa9iAC5FJ6j5sK8DTQW4AAwYzub5fk2+ifB9KyC
YVpp7lMKmIs6FmZCdi0s9zxhNq1fB0t89ibWlqCDKmPh4rQhF7Y0HI63+8YIXELJPkmIY3TvAKsS
KCpu1tUjdgKZffslDsLcgYuNEzkLcFgviEB14QYNRwiEFynZoXJAx9GqtHPyxNsmHC3S/FdwVmAk
ZrN1DqzRNz7UsW+0ULIz+YDWki9WEy4LpzU6HnD2TMp1DwQGnfQq+26Z/XGX2P/SDDC51PdenxbL
JzqeNTtz2e/8nZdtbX7uYMz6hYdZMf9FGD0o8edinFfMhtC4pNxGQ87MxzT+nNj50U8p3ALHSCu1
5g6/VtAQu/B5TWj/QEwAoId0YqHURJbnKhH3n9CV0ulqFXak9VW1K+A0deNARB658gDXI6EiWVeZ
c0uRX949f4tREFEkw7diN8ASVx2/P1RPi1xhyc5P6Oyxiqtt4G6nDpwCI/g462Nc8N4clvDqa35W
ndVPuk9fAufRKjdoCWHQAl0m4wioehppB+E4Yw3tfXWMVaEejlRFA05RIgS1aKygzakqT4sGIAim
/tS+d5vvR5Thi59fFJrOOyKQloaoFrTKWv701vpzRyQQqTQIOHdEXBLsDCyMM17acLIN7+Puv4rZ
1yjodXKcajGsS4iVfFxq1NRVP5KwUdSheXgYl0GTUfewQVdm+IF4KBZ3vf1nI0iMqeSSEWPhn3e0
MMsrWUgs5cOSQlyG2e6M0xbLFOUA4XsWOhINBdJqLCpaQn+Zzpy0oEzKXS9cGIRd9bONlXL26mUJ
KMquRSU9K1v7CRXwxcGfcFjE+VOnno3jtbwYClS3vFjEhXe3NVi7XmM01BLhMqPCshs3PXo1J8g8
tRRKqNF9qjFVU/Wuc5RLsW05PMga852HD4Ttyv//kaRQHVoO0Lg7SGUlkLjOFb1dXJjwLdDUuH8v
ZAmU5Pu5MLGv9IA+7uzVDjeHuM5SP0+LwFi+aLN9i6t/zAOllcim4RghXWLsT4zbcmxUQzwmt6br
q9klKfJqc2hQgNqPUNMrIs/jPSushFtAqEhsM7cj58iaRZBQlbvBpNDVA/LTINmEIB1+j8vsBeyE
hqgTXXJ4bP4b4719Vt0Q0lhUIwaxPzc4ebHbVb44kg/NOM2lqsjufHMgHCgEUdKS23MvmzwMhQS3
n1x4ZI3YyF8N07kocBzjz/18720X3UIvGO+3Fm2sQh9vUtHZoTtlsc1Q20Ag/j9b2cfA2pzyKXBL
6U/tH3jqZ1CcPHAiPe4IByeq5vm8gFdhg/l1/unA8UvGaFKJxjdMl2JSGgjc82GD3UPi0+HnG9Up
HJBUqTTqKRcEsnKLMrGNs32oPPbAXsDqu5zOx3jvCE26cOxOHqMjg791MRbHpJc1z/lqkP9DXWCC
0PqVUEyBqs5/MAcIk0YBqMru6hu3XwkS/+UldMyM3NOV1XGUSi5bvUayFsHarqdSWEIN4DheTehD
oyOuzOu6+sNUCSVXhXfl3sQFbOVo6UhNMifzBJhovphE9JDuo6H+zaTMSnh6eF63tkbe9obru2sN
Cs//JIrPtcogv6M2qMzMXrx10CIJQiZuPjmLiVIEDBdpNg5mg4k67dbkDO021swRFOx3yyzfmWK+
txCLt7DFJrQEImACLmPfuqlI6sWuICwQJfBdJuxnKr36ioVvh5MAPR7rIDunSgYeNmaTvNRXF9ks
Yq9GnSv5tYcuVo6T2tAQhe+vifo5bdcG2tpPcuN3aVu2FfFjs7StoPglagR+zQv7C8c+FU+73fsj
R5QbHUzGYWiKd4Ju+enZfYtrqHQ3PJ74n4d+1BjgoetYSL7Hu0anwmxs738tvcuCr5DLNGrz0ehz
CpHKJmn9N/R07E8LfrnbMBD7QoL5i7e8xzYnWhtNywqOWvgFnH8pBr6VWrrz7fi8lEXWdR/Ch81B
SDHHYhudtRe61UYXvgO2tTptFljcbbVaoP1haYNn0WAM7GPzOuvsdo78b4E7eTBwBBVhlkNv+30W
BRrz9rk4Sm4kOvCGdBJpRZ0n8U58IaBuPYDmR3SSPoTC6jcelJGya3BvKCcPTjPp9VWSK6BExIPn
ZVSGqyAUkCrkV6PenlUzXS6/pvf+rZ1VErjktD3dgVlZgt/s1LcNpa6N7GnDU4fOJUXM3XNGGnEd
ZRS6Of/jzUGKdbXdQeWS8r6FJrQH7Rn8HfQcbc25i9A2aAYat45XIp+0nuvqDQdM/xcvop4CSDsA
NcN2DaYT95N+Q11fOv44WyZBi1Gz4mYxNWOoz5WMnDs9T40oFKTbINcUhUJZVgS15ZuEO3o41bAk
GHEZ+bgpC3/hsrnh85ik5OXtu/L1Zbq+waSaHt+Z/ShZzZx/cpmysmV13cLh22TZ1bh+dJaBST5L
1HxnqJSI4V+Oh4vEnXW0cQrsODPHmqjiXiBYMaWu7UTBx+gwhBtSSNeJlo8TyLXh2CtNWsNrR44t
xjC+y400rE+j8Y6cvvdW+qdpc+yfKG4fLZfKSO7LZ7ow1n5Qdwi/qQRJvwROi5soKBCKbr5ArVvo
Tmll6819CmCGsIOuF7Cl8hvND4Up4Mx5e2YioyR6tU0ufMcWe5/+XaWOQw0kA/w08nBFyAwtn9lG
wBcQGW4BvdZ49goYHCKNgXrD4M3NNqJmtk6omVa+DzZmhz32pQxjFO4qRGUzD5i7Jvus3Cf5zBOa
AM8EwnJlJgeuGmIwfNnzxaf8a8Zi9WJY1YLBWpIECeVJ8vG4X05VKU7ce6hYBEdlTOIxAPxN8Xh8
N+RdD6fD6cSL9euOBLv34VNPoCkbNeZpwgI8tFWgYxri71Xl0P840vZ9VGBOPbuoXws2a0vN9nSb
jidZE+oSXykgubZ8FPrAlMPVSo+oPuyUbeD/CNxdqTrq6J38IxyGdzZ3ewT6X684Sf/yU50+2Eqg
uo6P1FPj+f2AA1rAnZYnMXVZMV5+lS3VGH5vM3CtOZNcPJmTG0wXcuXB6JMXh00jzFPBBB0GUfGe
uPQ4MLZ+Qlr8FpmzkZSkRQ5WfdcAftOp/arOxfqdPXhgKmEIV0kbuBWiEc40YrnfMiOLGsn2a8pW
uM44TpC24eYfDn+4CKawbnHrURzoz8F3Pa3xF3ORfvprvi/6Uc8tuikf9xtQal9gsXlSdp0JzRLX
idn3MgXUPWG2DNLWMEKqIVh6KP6vSi7dYuf8RjOS2SY8ZctZ1RjZQQlsXosAl95DC14exRU15yHN
F1IWK+xs6fe7yv/b4+Uz2Wfpxn0lG/F4WNgLYpfOgImfx6cjHxr2UVnHSo8Djc6u7lqnJlTfJyg+
DBJhNwcLMs/dDx7TCLMryLPMqpBNpRxfo2iwEljNYcsOK+mhbNuPrYRDlSiNMSSFremSlqLNhFl0
IkpHDDi/Gf3rZEctoJJA110IemwoA3xmBcIJLmk5x4l0rSLumiz2hpYXlrT7UmQqTjEBWPaFW6tz
8AvbhXQkpnJX4dJJ9T8YdZgjXEQLKMt+zCXhVq4B1C8sS5wcPukpY5Yi5FWKKYjO5m1/CR1/7oi0
hnkX1xcS81Aqx3kV9s+2PJzcaJ2b+xzZsa0NjaNPl9zPtLsSS26/trUU6c3nBYJr7LXYEGt6o1tj
H1RJyE3kYanp1QeQAjyXfVJUlrVbQmFuQ9h+u9D8VdXA+whRHztKTSIlJyHPOklPPanQg64FtP9/
HY2cjpiRiIVxYSBmuFI+nXtHbhH8Os7x+K4ht2gB9gKQqjioaaov4i0XTv8GCSQOhqcpgwKa81p4
xrjWNF6FWBpUD86tFA+58Jj1UHyIFNNgD9Tm3swSBWQQ4E2U3WglT1CXAFDx8MYtGPd33FwlGBli
vde6LyuupHeh00KQGC2wABjxVQmtX1tZ1ov1K3z5G9NxOKUvGRW0RtYDt36hXt8DiWKSxCEpBYd5
y0ClQMGqNUpFvwwGNjvvjeATcLT3MsJatPl7wgftAvLFv+Ib64wKmGz6793gf13c/b1mdoYy4CVG
QhBvBBkvTYQnvWQh5xNjof/MP4vq6Ykkvwio/Vjg9rQyLXBqNaJl/jHfH9BCdryAF8Q9tPay2nzb
F4/i4GdBYzDS0oxoHCwsSwKwRN+Vzh63clHDVrpN59iwkfsyohSHwtEa2waNNBSMBODHYSZGFpie
Ug69RkW+GyTfjuiXY/9xDuikClOGnperodAODR8M8Fp+l+LaJ+UiZu6ACLTvChXIkCgTieo8yFVc
a+HvSmVD5JgwesZULJTJDgrFASNLDDbfHEjIw3P6eh/TSE98O6iLe26h3/vmai1LuPWwrOoVvCeW
UP+sFXB9YZ8nU47FS/7ylL5qIVOzv0RCpbDHM4O5MImqdxt/zz57w5TJhLt7Oo68xebe2ls7stY2
OI1vAG/I87uuukQ0FQNeAS432KsHepIQVGnXexI1UoPIeXCIhllOqNY4cSUQmQ7ic0NG0tz3y0vu
OhdKqiz24Ypz7MIHe0CedqDQ5+z6ZHu2QCcpb+E3aIhzgyg6cdIheRtr+FdUt5uyXNEgcP4yy1k8
dpjrGKc9jvGHWu7VtOK0HuYHwFW8jDkiblTL4rDpBJNwsrBZEz/BaX5JqIsoLBJPy904ooxAnEMx
+WeAS952wgSTZeo6++YMg/lDZBnYHYltuPf+PiKGvLsm3Dw7UD3Ygu+YIQOAR+MtwhAhgQMLjKrd
n/JkVyYqydRj6T0JuVA0/vLzXVWfgJwKnRyty91ja4+S8nK0JnR3r4Tx1HULNd/MyJXhibfmLL6v
EhP74ouRbaq6rWn2KsrGllbznWS0/1uT7cwzqR2xlVZ9+RgYgn6dIQHrqHvXJL4x8TNbUNHnLhr1
AJLRAbUHBPg4fR1GFHzaSRjbC1KuVyVf/N9DFgm3CQrzEZvJt16lTuGpzUCfodzH/5bGaPGX1HDV
qtCMK+68Z7l6FXrz1T5aUzvneD81KT3LPJp29hXUCsLCZhlSC6hBKmXqCa1UVBLhR6o6JmhRZtJv
93l9JvxHwfX+AekeAKQTQ5CfbIXzCW2YIa5dX9in2f1SwRDi50PW6QgXNUqhS7ototfxLkewYfEb
aBmGrDH9F7n1i5Asp3/VbXhjHm/OZN0chg0LULGCxB/crnbidCalBHtkzq6wMNX4Y2z0tJukCSmc
9cPB4wnChk3AST64IUP3InqEwt58FNi3R9fCwXq4rkhQhZAvRhW07a2nVGXTkzp09RY6pMXf3BFF
jf2sHqkIqRJQTxUZdSiki9eKPw36DdxlgTMvZ8MIO35U2hWa9TbuPFWwhnLIUdWLgjBwLZMdjiOC
6iHsDvOenrHc3XgNF8wPVKHxU4KrKUn+TK7EJs0ma3I1WPnaObm7fpY1E0G55Sk20BFQLNI6hyJV
Q/cKnsh7OGuvo9frrizwItjv5M2nKBxoLdyDSItpgR9US4jYTKjESQ7+w1btjB2KsevYqY3b+gZi
xKmmapx3jZQnSucafuN2/IV3A/7+MA2R91Zkypw2lG6tGAUrT684JbCdMv2CYpHENHfUAT1IdO0/
ODkRdPP4/nVTgnL+3GDOPJ1E5slHs8P25xR4Gu8OtBNnQrtekj2FE904yho0FKzGisim3nfZDhOf
K49vsR51d/wF1YFk/s9mzX64BYb7984lvrNq1I0U/uW1N34rPS9iy59o9oFqI/TpFxxjUMAGumfZ
ng/mOEK1QONwgC11NXffQbwzn0IV3T908a1CRPWADiKuYMUgFYJAAOTR3+KJ9tCAybMWMHvjc5H5
uFkUPaiTOshYde5k3BuY2LPuo3k6ijZFjffYaSV9cV8WK6Z6/u1R11hq6sIatmijteEPgaggVDvE
BHNlKiHb/K0zrdBmKaRTwWeZpnMvo5yAIJj1EspyUz8E2/DSezjNbzIDsLI9vdatZSA5yggbiHx9
9G5LayCoE2oSzz3BlJB5PmVn7lSFKaqZzuOYxxyqVMh3cz5XdMP412rxbvyeDRcOAeL9c/DWft+1
eyB9v2MPc+hQ2EEgK0TSjkcMF90/bSjThFk+nprTPU+Ah8JkHMeK4plZzlLi6CK/FNmuD3u3i/Ob
W2LmXHV3TPrKyC+8i30NnmRA0CC2ZEduo0SYHV+lpoQ+W0g1ySHx5Expzfm9BuRnmcsDybOzWBar
jYpwfb43Pge7bP3mtuZAYuAT3YhtLDDQF/Rn+7mEdpcNBmC++boOrrY2EYd/e7HTBbgoHnEqgI/C
lmgfrjqIMTyNs2LHbEO4fEobNXuUjlwDOU7H4aNaXq5y6X1kYqkfBVIfZDD+BkfAntHeJvo68nBc
gsUkipa18DeTivvx67sMpu2she2ou8bBR2mve8wqCzP3WIffVgVkyEgiMzcH5ISfBlqH4Z84cSfg
ioYrpKor6Wg3g6ZY0/EXoAxzfn9gUIoQtWCGjMOlovQuaAVQ8D5wj3e1hqgKDFJ1ofBNaOU0cot4
XxjW7fnZ5P4g+l++p0f3OSfEw7MZM2C8LrrM94dgmGk+aq805+BsoL4JSsjWGMzRgPP5Ai1TstuG
bWvnxWaEfqU5HapkM8fdaT4DSMKsPWRI+TWBxEU82nS6yxnpeWkhR4Zt4luYN9y46bA3ZcCzEk1B
m/slrRBmAcvO6cGnT6gZ1ClIef5uTwkNWGW/nTMO2Di9laatcylJd4HWyFsKVvHUPUf0/hKCLzHV
+3dD4NuHmim6v0ssLwTsgQ/rCOc9P+9iC8SHpPESL3uFpXe58vx0CEebTHvWA+j9+9yArYozvqla
tY59IfbhdiEFactJuajB8mfDRpJCUYm0YCVfvuGdq6MH31lFdsNmHxMWDpnKAEiZhrUAgfuRbsKO
/8IKTG7EXgNpy7TD0Xndz1r14PeZm0lazUvscNQP0fE6CN2BC6nCHVc6dgRVmSHbLZEQ05IHmCnj
BUE+npjqMF208mGCk29qsiWAFS9pWoy6FJpGp6k7NbuSAXYUejKOO2LwUB5+I4O8r0+xoMlk7M1y
9/KbS5Xsnq8rJXIauidpUppThJuzCNFPMf5kQOWDPA+n/iD/+mZPpFxD2rOiM5pCe9v4hE4yIavJ
RQrSDcanTmu+jqf40KpvnSfIk4VXrgSzPTgp62Ergsa6Lj+XlvgQD765qOB4gT0b43evWhsCwQVI
0FIpYeGTD042uTxndpgigHzNzsyYJLi6I1WmSJEqmx5D93WyokOgjnCS4ZcontKbQ/5sPLFsSOha
RdQTK2oEg7SCcUbt1IBCmjsGFtFSLJtR39DR0fTjnnw2WEROfA0gvNvqqxVWdvhwXyedcQ5PSWZf
8SIGNKx4lcjBX7VvXulrDdV5OBDrYD6T/h0e1A06mC58M9tkE8rhCPze8K9byGiBKflmlv3sepDd
/UTkMItdYAAwdgFXvn0sIreotO29Fp3YAxo8D8fr388nlakMbLDzk1yyVU2IHOMrRcTV5CIcHTAV
G80AaTdsBBcu4I5RLH8NwXVsG21T0rFPLbRObtwwzDp+rXMxXBJ4nxLs9jDHhhlaxLDpSkdLUhw6
aua1hiSdKgCBH4BIS9bLnnc88siZdyZuYXMqPIvbbWlXJCwUGxhiE+6kQLsGnZw+BuVEXPoVLcte
iziKwik1hmFQWGr3gMTSxgT865Z91kWXTPvaXI6F8aLzauGuqiL3ZM/lHCaRn3GJF1LE7NO7zANx
1oSRloL2HPvQjFLyxHwm55wq/lJbeNC+T9PE6fyo+N3utL32VKPHKUTcYmluV/zWFud3gM2ya/T3
OANx7lBQRiwvs/c58GuYGfdOCxCA4jvQfEn524tHr76BFjosQiF/M0LLtAk/8CWgOII9P2D5gbs7
eSjiDnTboh+RU0Vro1Mw+zdZpA/GPKTrlEz8xTk3IczthCDT3WWlcKm1XxPHu0j+qmL6VA5SJFOv
oZsff/kr5eDgdyFuY6WKcdyFh3/nAz8nGebmt0XM0lKTMYfMgE+LCAUfZbKFTB5o3UQDWxGP47Eh
grOOiXI4kRRe5ZCb51jry6F9mOkvnP/7RMXNrayKLSxvvfdqbfjBMWlXCh0g9ZJSgPsFj0P+nAaC
61zaoZESKmxYQvBZrU6+VBvbhpb3xJ3DJHA/1a9vxGuaiZgnJ/0rPiyDMiemU2HmwFtiF8HTG5b2
kDzQLpLqmKsX7U1jmT+660g2fDkFgIfN980JIQozrTFSJypfIUDAVU53KoeLLONOQbnQynyO1Zf3
LJt9iV5H08Bsi39u4mMwlSyqMk8ABfBSVF/Qusoc15wlq9B1M5C19EwXh7ivWre7fR0FFWv3Pw2+
lvoi37xC8sMbtZyv53qHhKuI+rZmUJ7h+55DXkWk1Op98/WaN4uUr/n5tBkY8mNsd0VGwZl6rokW
WbSHk+RUwfuO3Sw8F7Jeub9bIStgHI/YLWnoYlpElV9X1acUTNGJcWej1d2IAyydDSnHakmfj7sa
tNz8mYfkG21hctDZjyzHi1Fk0rNR5OyRDRnYq2sghYpoBMpXgwGbAe0Vf4C1dwZiiHp4SSlm8xAL
EplXn9HzTGXmwuqR7aiS4bbda+gCRPSoGvn9UL1lSYQpyTKVhGCd4a98rXp8XveZ2AtKzF9CyDWh
/yvU0HtnRmmBnjhAHMgPXz+AsxwY3hvkEkd5KsUJZZGi+hlOH7K60rSZU3Z3CIn09SPjBgreh28K
p8uVOkQ6k4I2IJGdtzo9O2gqqbJ11n0gqfUcoY04qhW22V44AxVHAMHcx9jcXuPf07aUrvpXwDtV
2qWU+emq7IFcwkzr7Q6dnIVBVG0XEEMD6P7m8NHdQIgV8nhBqvocK6XVAW1lNEGsWwMcFZ4Bfgob
rftLtnb4Tncrpz5j4JcubrI5QhWHzmrZyljXKNoF/p+yGg24tdJTsCHe+pRA3nRfcGQMMk7gH2kW
xrI8Jx0XprHA6DxBFA0FcmtAawUMFX+nmXxkDOdhawYgIbwliTP2lyCrUhI4k7WrzE8cCoCRJL05
aVfvCazyNGFyZdL9ufyMqjB7gH5OrTRQxrRsTLozSQ0WxPXvo+5hv2wycdoLEDyJRHVcfI+NghuZ
S/NSGWseanf8a9lTn8QrxO5eZ7sSrr4VVQ6kc+Cd3bZdK79oTPXEKUCh9/LyDqb8C0Ib0mERw0Co
ZESG+cvN5vdkAljC51ROSJMYn3/UPpRO13MvShwwtZ44jEK05tXFP4R9HNYANzPJWCQK9fjARyjE
FAB0VutmLglyIiqDR1kMNEuxlZPSevjoKMRVhEexUlYcowSBWPESVKWph9R6LM8J640+4BaaRvfW
wiF/3u92/LdBTAasY3Yl/48AXT4qGvtOS4fCvKOJDBAO/VKeUTXeG4/N4QiL5mFbM0H7z921Cdg2
/hZPJKXV9+nY/6eKhxXJp2EgBlX1xs3kZRY3TMazzva34VVJEGCL0l80Nk+iJWctfvI2tchkeylu
kJP9onbedvTzIYQP1W6ErkUhlfjXHOWsczAalYdHhEd0XV46AYpY8ryo+iR9kgW4ebjgv7GZ7OAi
N82se3Xkrmypwp5zc2bqMfarfZ/IRk5+ZgCOAoIB/nB9hfgdLLdKeObffr3Mj/GnxSp8xpT7w29g
fYdGH+j4EPgKA3ckHLLZlgH0vS+GL3g3LIAkQRAY+IIA0n5LH6P5XXtaDuojtHmhpimtHhdyKct9
monvRA4NKvlzeDuBalMFTwFeTebC+g9NnAft0AOf0UHLEDvm1rI37Tgm75Frt0OxpVr0OCeR/1MH
ARBTxORPDz679CIX4WE1QpES3Ctj8SK44Kn46CC8LT2ZbIkJJZWyGT2rga4ltRRs9YgoyqpzGl4h
+XpsdnqCmwQdNvvBZ0RCKa30JJCezxxWTxpJRO7ZMzNAGy/V4d+1oRwwMrGYVVKKjTFNdNAFUbg0
d0IjSvCz3gjZoST83DnV0f+rdmvyjdTQ8LgT+Ay8MHtwvrZVUryFTEz31PPAnXAm2WJBVzZnf5vh
XEQD7PLLsYN/WULp1i/FPp1Ag5WmNAySSo6CrjOGl7xbYc+vt4IDbHwWtq7iRm6VMaooxz/fY33p
qdrNhbdFJ3aUDcJwqMnLJe4PkZM48pFyzGtB5/5pG4KEuj/kdhvQg6JEhN3z3Z5vRrHoxjHC9ACy
oxm6mXlLDPIIj4McrE+tIafstygmrZMjuHIWxwF3PVUwW/BwLgI1FjPixBaSs56P+aSGy5nd0Dhj
EHGR6ZX0HDJEujKWVMHgcZGjUobL6myMAyu/ib9J8+OaansyBqpB+Y5IDTBsWJSTydfRx6vxsPSL
AaXtDRemecdotVqIN3QQs0otdD6tEKkeazwMp9TLOtriljWFQNWTauQPt8/NJvVLEIvloJJv464T
OHF4d9ExMasflgN+hmLA3MTSwAsv6aZkF93sfD4aGN9kREgKsK/qOW6h4Sf+u8UrbXkRnCCywi33
QIMwRTVamr3NO19Xr/5kcHdU6cvmZFRRoMmOqcDRydJYBL5DCBjWPUZNQsL9XwvRGm/Gah+EQrVC
KYUsfnHwF8HDw7l6X3fjux7ypd4AKFw9cjwb6ZHqWmungWh+1eZJVPqwwQtkoLl7ctXwFsbEbUQC
tiqYW5aRNYmYambf6fJvNI4tgIwkyUWlJtRrKH4hcc5UQrNthBMNBhPxoPjXnxz5Qpty0y1Eo2fz
Jten3YAhq7kWb5otcH6Tev8FinzuXAZHjWGpsgXhSyPvVL7btH11upOSy5QiigNDtwE5zPZvyH2J
oU3h/9I4cK/6F3NZ1l52cBaFmvdq1rznwb70IdNzbwYeVvNc9aCKqgED/euPn2zRQiFkui08W1WG
DGEASAUi7labC8SYRnDzWDf1RUWWUmP2QJilcGPLzSrfB81opoZZFbspQ9cPLHQwng/8NIa7iCX7
ttyrqxp1Q2KEr6T794+/UI4jGyfxuIdE1m03WSS9eBra5B2DgOUB8BUlncq4Tqm0CgqwuGvVwwuT
jtTdI0wI8X0ArnI2hVSLBLqPZsZzzqS4Hwj81zoVSUGdJWZlgsjPBRtua6SOOSJ3kRdTUG9U2+Kp
WJHJHvPupg3cERUQhDWXwbU41WKy6uHgGIEUyKZUfYIn1wo/3uxLaEvHKmp2eYYh2ujsXMF9Xfmm
bCIN/58E9BemLTtk1XMhjcFQg8JJnZODw/gUS0juWgiYLMe/auBS0QOtHgRgy7RRG4YSQatwj7k8
S4XuLT6IPmluHts+t8QN0sr2XPaX4ccww6qbU7p2pCxe9fi7rWyiAWEeA9NpB993TEV9q91GGwyl
3NVIG5atMd9VKyDdBczffSJskLeAg6KEDuA/SJ2sn9cPpsLEGfFJflwemz/N93hcuIq9r4sXa897
FNWleANcLSlRZnuPPYQMPOExP1l7MzcDKd5LBBRu94gcCZdkrnrlHO6dmrPal7G+De4wKsxe8MPJ
JggVv2Kmm84cUkYjeEVXYpf3jriBbNAA6mSJri6TDNVxxdWVqRYqRs4VQWIDZTX+T6c6dEwLPVeO
b/GcZQkuHBwiflDeN6TI9DBTZuJQwnBEX2+lA3cELzD0y8euBArjep2Npc5R5FRzkJgCeLPUiZfh
bN5ANG7gyUH/1R5npQlq31OvxUcUKge0l+d73LvMpdE1yfaVS9AGEN6LqxG0LLbPmGbDrfPG8q7+
1u27bT21kLIDbN4cz16BtzJ5Xew/m1StvSE2bqX/hZOSofqOJMVS9BD0SaIvDQ7aUUBbSg4clsdy
v06XjlnSccAb0HoNGUSSe7+oI20/9RVl/FD7yFdsE4H4T3fd6ftQ5JmyM5ZLD3Ct33pFqZuq/oIq
cQiqsak7DBCsSJaXHK5bHq0vumVaQ9qs3xF65qb9rpwmgmnSLDSaae7zEzJdTNRB9GJPE+t2mFRN
BNN0C6Jh4OFrP+jzzyFUHpinHnbRqxCtrqsLxeAR6wqTbZetfTUeSDftxjbuvyV8DdJhYFxPG2Y6
UkmQ/wH0RNMB66FctXN2+EmJuuby60jPbpPCoSSIZ18olUeiifFYwImr7a0g8snzxyvZBd5s3U5I
7Hd9C39oxqtYW/+0WuSo0tOgSMv/V1EvK7SS3YM7AgXA8pxZZt/X4FVBagsxodZd0zjVQhQ7rddE
o6HpLh6x+rNRxzzhQo8RaUIvZnkOaMHfoSx62MQRlszJc7phMGjBUcaqeWso6yz/3O9AZrdh5bDi
Rpps+INV4Y5QnoOAkux4TzCvN/wtntml75ZhhhjTOr6YmfLecT3KZgElcd3yESM7v1nbz10rfauR
xhOwv5jgNel87eFKbTDpYoekT4D6c8j2NijZGkFraxPdEdYqoYqUqFmiTQC8S3jfvMrwNXxl0a/Y
xZ44/p16RaohLIci6WjVB6ySbxhE1lr9l95jxpfDfzTMGRvk5HBf5MySJs1tsYP5JVc12vpEDeMO
YK7wBNPjzsXv9j6aRw/7Ljud7jyBc3XpwoTAto6ojZaznUGni/OsMEXRVn2l976Q/SViNA3mAPrF
OxZJQJplsfhMIoRWECHkYh21Gr1gItfW8a6g96RHWCo/xtzyGXmFHiK8Jdo+14Tnj1px2zF6GXaJ
YqXhZ4Lj1haIDH/95fAwWIdtOKA1SpjVN6OKwANF8xEqPl8CdKT/50I3ujoZSfjxg0pxKLcJZCvo
P9+Onk5m/wBxhCSb9cIthO0p4F1n94m2FboSxn2qyhp9Ioo2gXVZ61W2ecDdDj7Q5yYNVtoK+ED0
0Ebf1NloE/EfRSQ92QHD6wyMjbealGabwy5uKdBmpRa08xJfVvvSsB6dXq8bbSHbuNbf3uXi7ku+
zLzX6WByB2xTj5hZPMcTBrB+n6+hpk94vd/j9z3fY0mIhQfsKGVxQrpC69Qe5bJAZZsX4x2EvGDJ
kFsJV8zSXEbmdblZDlN0RpMOfoXkXn/esm06fbH2R3Y+9y9sQJsnv1wHasEYiA+3H1y2XONXu3RY
f0EsOiLAZrv00cx0d0PGRlKY4DDL02tUTPHm+CDwwZyQa3FpKPxX0V8YN3HycBWFVxb3DuWBmY82
soJIEviyEBa711qdQQ2xcuIy+ZjePfnoMArWY7fU7DJhAy8IyUZtlZ/5LiWlN8gsZzunjEeUlm9i
ObRECWknVUNQ26qc5g+dL5/z49QU9LEzjM4hHXllQjOKCfNdSP94KeEMygJDjXQVCmMZhJJrNFoO
76XTx+smjWAyzBTZCvTLlybLvjP1HWdYEfRlTeflaUea7NWE6bPcLx/CHcg/d2dcmfOWBK/rXTNq
Nk4C7ikaMn6NkFFcIO0mX4x5m+QYzYDZ1wLQCKAEHgWByN6CNELlnPD06viVC9re65c5zSQvcYTO
a5/B0Rcki2zxEWca61Cc4krw3Aa0fQqsxcTDGiTzTVsevOuM2l6S7AXurO/K9Lfa954IwpUIml0u
M6s7Vkc3K+SANXedKPxX52Lnx0EbI2BbfoKwMfeIYZIRPZqTopEJKX3l2NfdCzXuTHkPj3yntHx4
309oOM4LcnRg6UOG4P62zkE9Vm8a9aBGsx91NFl96bDyvWT9t7zaliMwAgB5lf/6WrzDbT1WiqXS
Mv0q2oul3zsYq/xacPfArsS9rdZd3Mwuskx+wfbnnmPNiVz74hfqQcTTQafQLaW81duGfCQac6RT
M/mdacUwisFUF7wRH7X26Z5QGMutirMa09Qc+KrPSC3hzreAeLKyCvzcLDX8f3moUOT5J09DHLs/
q2RgLP82NP24T4NSDoS7CJprSNKvV7Fi718j9CMICuQlkUy0qD55ZLy6bCv3AyTXTT4LJXpFt8iD
LEHBXYZMn3fK0o+LEMVJAO8A2CDMyPk8TMSLd/RUo/nPPTbPtEIMNffiqECiNhMcxJFoVxBuIT8c
Qjs5+532yhMg1I+pDxjJst4G6nFVyhdmr2JbrCxtvMZCca9Ex5lbyg4jkMfgXCQtW/U+L69+qBI3
hGMa+D0ivUnWyBEZHPT8WSPUTcmh6b43jorYgY6IAAMM2TNlElOlxRNUgZx4tcdcyHEFHuP80Byl
Tf5bzhE3T6LkRD2i65Xm9iIGDf5ZXzEJbvihJKxHctE21fnN0zdCWB3KO6N10XoWwED/vLteVHu5
pGbiCjk5gnszJ1G46PlDLANz3sUSR2a27WlqO3B1mc437XyAEo2lB9HD3YkelJ9NCsqn4nDEOUNi
4ZWfQMFz0g1N42JNKFhWNEbMk5TF2T0w8S1oyCh0Ev7FFuTTmhnZWirSTFxyIkQwz8QoD+fFmXBi
MSZnr0sSQXyt38pWSvic/0ci/reI0s+DVIbONkmEPGZEV90vXPo61EmLTQBccBCMWQub2utTTpfs
5Z783IckGTCKHZUScqmlcnu5oEtCbbdz4YgBC4KpD+nPRnYgy/ytnIEZbIfEPMczieE+v9B4sHzj
jRra3LpvgYfZvg4bQMBwh4GUZ60lm65WHFdk3FrzUHt4ohLYFvNC1YpxO2fJ/j7Y95AD+cbfhOHg
Y9bq2sctsOxT1U6MdJoLhpEfTmNgn6rlmwiJpCeqK0e6C/KAnogfvQOEnw/Ioz50zs/UN37T2EWH
RIZJNVmJXQYdFHVO3kPIBAV76/cykaVYXZ/P43IIGGROfJgF/xJ/qsrI7ucri4rNJCgifsC6WNNZ
MHjMRda9eTb2/J+iL3dQx002c9z1l46BwxyfJh9tlnd59i8bOIR7r1uMv+IzdaWNTM/ZEtEcEuhv
uaXdtBvG3LJ9Y+6wIs+L+dj5Ayyxn+bnZGgps2W/quBgxoXozLavI41Vm3+M1Fdf/5UJ6eNbYdp9
HHRv0Ht1wfvS2CZYOQcRxquJS5MF4FFCp8GyYl1zsTOEO5+n01fLXXpsTfjQcwx8eBvTwhLBxmnb
upSuz38Ni4etAUgUccBNRcBu+Gk/qnvrt9ZliqiFbIuTZSzw5RGHlVuF0NL/vadyRb4uSyWke6p1
KgZ4TtshxtFX12xCH/dCfirpnnrqyus44NMZYx4BOmCL0haW2wV/tNlyo0g8VsVzN7IoHVe1jFpd
i+tjZ5uHVUSdB8kPT+F8sb392EX/xZSXdlBGOm142q2fLE93hh6bnlzg8g11YgMGwzeKgWEN+LUQ
QCLZY/wsApmW93TLV56QKnKKA1eyL0vIUzVuJfRiHuN1UshM2P1cA/3nHSnXS9+q+R/M07jwuAPP
ElaRPUxlFoyIDupvej36qy6o4zNH9VDIyNvRSNrYDQEplySrOJD6Sl7MvfNr0fyfy/I86wPpCV2Z
F2ZI7G6+cFsjRt3/uoQxT4kyfg+xL/HNAVRioIwK1NK1ykNjiLV++GZBjmth8CCPjVq/c4dr/jN6
JDjLHMpzFXw5q3IFznnROe8D4PbmFTlXVlLqvx4vqKBJ3KlDAkfpl4gtySMEP1xExkF6UVtXe8Sx
dczLamPZ49GTJNz7Xvf9gTJvykmgJVoO+GgvbUZTJDuzhrrDsoW67HDcTemH2eaNWx4396MUSbdM
qEoA/CdDcTRYYJP1wVl4Y9azqN/KMoZEnim0qfHvj5GJkGSzxt0E3Wq4ENZu2DdcpgDZS+2bmC9h
DQv//rQB5buLcvCq8UDBEQN0xVF/fenrJQQOES3GGRI5xrXFCHyeTVF/jYcK/AncLu5LX7Uia3PP
xRDpA+UUE19LKLLWg8lKJ2R319IMxVXxKn93MD3i0kG5J7+nQD0ZbChaxq/ZoIGaWIPLbrTfhxok
z+BQhjGRwtRumRq7Tbmbj+2rftaTxp7Xgvij3R4wErICuGRiI4dZq7aloybTbe4YREuAZgEbTR7y
irh+1P5tTcVZf8yl5N/TrCyrlaunnIvfnExs425+vJHHchoEsuhHblN/iPt/Ib2RI4gdbXoa41h7
bQ8mzcqfo96tqIV/XCxFCj3gQdAbo1WmfiZ7NQb1D+KRL4141V4nTdX8c650LvFgp/DPuZUKRoMe
K51CGYSOyYLzoHQhtfcqJW7CCi24pwGuxBUgzt4YOIr+/kpLXNNKHQ0j2MAg6bJ1YjcGqLDV9iS3
jKnZIoIR0gHUfZpbT1Y95YS4PVKAo60c7D18X6f4hgh1+usupm2lq1riEm+yPBAQLKBNIDJr2fST
CjzeWq8lTffbBVQdtsYuvHFsaRK1LJQ9fGDbptA7sEvefGjvxLiSFp2hobfyTWXgKYLh8d3r+QIF
TFE/Ji+LLnAxUnsb5TNu2zFL4bVchZkySi4yfcA1InB7gfDwddVoZ6aO7J/1aXWuF4xM4Mg5+xfY
c5vvBT7Xqyy8mFD2xXUELJdOeQXfK9KhwGFCNqStrgkyXyv92sXdxw3P3GZAL8zK3IlqeHOGLcgg
PXPLf8LSpypDQZcOlgdR092iYhYuyu94fgY3r/6vsovPDfES5SFutHGDyuTu+cBhbgQCdaUgmlNM
ChMe+TfssPwZC29dIFN+mblHtZ0gUXKPum1uy+waLiwEAlUeahJCTqAa/MaIRNoyzTSRXeqtu3bV
QDdr0n9OH4o7ARU51RdkV6tQPLRaWNn/qc8xg7VjbMeo8MysgWXwzAuaiTWh9WOOL4LMyk4NPizs
LKOCahIHLk2wh/P1cPJ0evToDx8awtb9gOw7kSwunUAjwVnvsDamch4fZAKn4iCUmR/IABkSo5O2
3plbqQ4LIxjsuB0UIB0nhFLIoiONpn1X0ADLe7pnlt6jg34T+yhE75PASrMdPo0roncjmB/68f8Y
zppxOkr3dooTgWr5osaSawUw+VEIIZYE5Ro95THRn1oJBAe3gmH2vfL1hErC0mSvDZv/6aFwVuoi
P0wYXMkW54L3o2TWeLIf85Uc5DSEobA7HKSf7J1CmkG1Y2z3fePAv3zaXFcblA4AmQ948v4aalO+
zzW0a3PSPbeud0Fl2IWj91nPoKv/8ft6cR6xHXi76991X0gYldI6wwbu/6/Rc0+0L9sWlMXc0+WH
5P/EcDcYDk8LWfI7BkQyxYS7AZf7gjEcB1Tf7mEAz7IUn7C1o9Tdc7loLQgtS++Y3NTTWEY3suuG
Yi4kYV4XtpNWhNGyb2LBET7GLzSTL13aLVTP/GqF2oroKPI/EkZK+OwLKztNYZkaHGbDlP5yM85H
4lbNHuw8JC28Jue4HpIzviteePd1PzxHFsztCZ+sZfksk9Q272Fz38YuarviBdOjF89UsdrhdoDC
5bfykGbi21qsIHlGzUGt1RafcxeIa6XPJXtVAJA4Ea40lFr/g6iV0cExF90ALDnjziCMmaFaS/20
Nu60/7oGXM9mjW6CpDu/OV+N148gVMvs30MDXaskgQqm+zVJk0A5e4usxVuA+ElcafzqdEWaDkED
vDbLP8zRLjGkBBUW2bAAR9nfeFcOttQEBLrYoV+84yJlGVjkgmrOBM3qK/Zrr5I1RqGO46Lcf0/l
YAZ55Pn/H67FEIxMwAlyGGWafYu1B9/iWh+vUJvbsrb+k6eBghEPnhoZXwnxuyIHHF4DSh46bsdk
iEHbzCpiEaP8Af7OgXjQaT1dC5G7EApRRaHfhrNoYqe/ReyTbCJ+yyCtd4wrtQX09WCWMzurPFha
BGFBiuy3N2jogwvyL0z2W9DZfVmMsqoDuRn2cO+p7l0wV6UfpJi8fEmrSTBzyyp2rHY6W+D3EpWx
KAt/lYgi7JUASkSkx4w7xBZHwq9cegD34q/cHjTeOCS2ESnbtA61U/qR6g42Jr1ylHd+yoqO1sHW
VnMFb34FTKq0EVKPqRsnrwztl2JbNlJT0V5k+iR2naJiCkqJBmwqNJ0JVmaDoBZj+CKCWxgjlhYE
Nw2JRaacFEbgEwMJX1Z+uE+mGjF+gxEpSkbL/XAN9FrvufpsEWCbChJ0jw6Oy0RRktYtEJNg9rhR
DQGEG6+i+aObj1cKFB7Aab+XKbwR3Zm6NoE3ypZ1qaaV2/fFZZqaskQI8H1PGgANG4oS4bmkD3w4
C/lWh+yKzNwK64LoarsduDe0T25ZRHFTg6dODIhKD4bPU6N1IkSkBzuZYQ7eABTKNAZwVYkpPCsk
41smHv0na56fw1tsziuxbRsqUSBiEEsN/8PzeoWhohlV4HVYNFNy+HnmsM1PB7ZPQuW1io6+74Kp
SMmbetHjQlQbDQht/YvEileHKYW4mK7GE7by1XlywLL81z9+flEW3RJMixtIMbLUV8Vrb9FyD7tN
zU0PROzyHkx6DNskTZLhoetNXqnPG9dvvKYF8ZnbmCY7F50R7RLwwn/Dy8ZUZfrrTA2gtla1qurE
OwzXr1v7CbLED1agi2HuSS0WVxug9skT6ShuwlEul48NEmL0GQOH+jiAmLYrLdiIo146wR2go+D6
nuaGi0oosMBCtcAAelqa96gMQlQdw+kYXBnu24R9XxS8nMKQQEXMPLWAPCw/3Tew6SRoxiHeqvPR
fLGmRmxFYuMBqIB4hG/HgXXim+eGA6XTHUK+a8jLwM5GnjUQpPZmeK1x/MoHwzSnLcYD8+c/eVYy
uo/WnNXIxIZ6uQso5vsGWrdCIe6AYdND6w6cwlVYx2Byl6kp6rb5nzPZOEPWWLHv4jV5XoXGS8mH
Q0m6DFisWo1Td6aTGyT6j14/h9118w3maO/sURJkVhUz1qbpU9X2EncCTf9h8zJx88u/So+jN5Y+
5k5AEmRkb3t/nPknaRbxRaXjuj7MU7IjcryRkhiR37XvqoL94HHn0m5sdZ4P80n+YBOuKnTty6Yn
aBGbu4zYjsoLK0gwHV8x6abaoSCCMtkvgzMjtDECYZ5ytf1PpI5pbqoRVegQYkEsWcb0bfw9hnfR
PwosQ5170a6ZciEoh0inEwpHElJ1JVjNa5iHVhWrvXQVhTQI9+2Ik8jPs5FwdIRGn0VJDD3XG1C2
Sf8HUeKrlxuIMWHE72iGSWr00EBj2KzkRbhyzH0M1K9eKCzgxYJl+hF83EtxCt4oArd+M5/wUdKK
56YlZMtYJXDmwq52T3kZylIosG3KiRi4zld8mCy/Kjt/MTLKvvTuWeJ8ltGpD7AaBpC3kWo5+qcP
q3T+B/KrhPy/V0BgZw5SUNpnZ8CRxWbpOXr42qxU/778YyqZxyNKmA4kKU4/eryGzBFYMRvBb+wB
hAyoFYXEqlPqSVxL9RznTP5L6L15IruCwbbsGnjOVA0qbGHfPXJW8WnpCgpNfztCjCjOnc6WMoyf
r60U4cV0C7N4kITh5lwrCaLrn1BChbxPTkOJDcO20SSQIKYh1oH7U9Jghc8sGj6fWkDo5dn8KUne
EqqSmqKmWTg5DMLMFDVFn9oRPfcJ+p/6z0zDCdxNQnFNbfSj54/vtfyaD042qsCiNBgMMu0LV1NQ
jqJD0wVi74YrLaCRXlIDM3EcUuaXjO4ruMYZa0+b6fifGzxGLuQIcp2PACjnpwv8t23lh71qg2Hm
j9kZmCQF0MT+rZDxjfCFdrza3jQRfYCsB3UXpYSrLIh05n7BfnHhDc8RGmS5Y+v55H4eu2fnE4ql
H1kccwRouELYUE/rWCKmC424k4808LoV7toJeM01eSJmZjljqjXdZXsBOO238o2CTTIztdgOIHJE
PQYL9ZLMtwY9cK6Xqyxvejjm/hG7eQ5wLFP67N95iQe3dPOe5skwH1/nFU6epAJoZU3SRf3uSe//
+eTNhHnFhdcjG2ki/dfnlYjIrSWcEEu3Nk3cxXTMaHwGmpWJhG0Fb9XNXAgvL/MR85iiV1S86uqs
NS1yiMEk2WKzELC7FBdwWpoVowZRpS8lMmyVAze0XunFk/bPjgRJVTjqMjaYZuLJOrNGNR0OY4Wo
lct0a1fvhHzhUxHz6FUuFyteWnCRPktHUKjF55MbCfWey/snIzKtTb5gsTl/MvCHhB97mP77gjk4
xwbD/jauLYEFZWzPXuxI22VAdETnJIdcr+x4yx0nTmY2Fy3JPBw7ZEllvlYQrmC/qJ5y5j7APTJ/
CR6anMVaKT9xhNK/Rl7zxB7cFEulZ9JvgvhPzR5/TBdv6s1zZ3PiOPdQW9FxwyFUO3bX11Rg5CF6
OvQ/ct7GIS18QzXgwCELEax//3rRMmJkquKdE+0GDs78D75w7SVxGN+ZNgfyiSB0O9PG03D9oBjy
FaV0mxpl1xohMtqZU3Mdv2fXNG4agmPZg5GDR/IDPv5UqlMgpX/B4kYPM+XYT70kQEH+VwzpGH8j
E1PMJZ4a8kIe9RKe5ZcnlBeAQouFAl6WCAum//Gbbz9jleK92QuqSv6Fl6HukGOI1l+DHoZ2qr7H
hDJXFMXX4MPYqckvLEu32eUFnTzxuYkHQa6gtHj7xPnSFs1dSsX2EUtNdkk6LD6qHxTE7yk0InKX
K8bxjZkG6+SU+9JeivTWoOG8ai/mPx9dwVQNmVx/RDGm1WqCQ84DcEdm+VSRU4uj+8RaX9qrbVBf
1SxP3zEo+LdeL6EOruIZ43UOOaXGPQhgaU8vh0t2B2iQVTCVYN7b6Jq1slbkT/HxjswHal16EePe
o3y8fr0v9pLS2Uk4yENM0z0XOI2j+vUV9AYPCArhPhf7YfOgN+5g8iOM8eVaxKD3/s2L7PATvrka
0fKF4gVjmOkXftqkAJWCpr1fGje7rfeeZWeQPkDYUdaRKYaAdvUxGFNSXhWZpQA9ISnju3+zfk/z
6fDTfvghXMndy9nwiUasIJyWllE0kGy+e57cmqsYD7bKvJlFZzyEJs8EWGrEBFrjejlcjLjfg3L0
3F2ut2z45yH9b5FLTfZ1rAptbHFUF8aaJPee+HVh+gV525RMwdRdDhpnqYSkdMrAeqqpL9Si9Eps
XvvBBQwjyL50Yc7JHz+YQgn3Xo3m+q5I3bOo0Kwyj2cJc1MoKJoIwTnvLaxx2WRAIGH0zYm871uu
zIgwszhWEDFxlUYNLPncIh7u4nEbXHRR4A3PnmNortapTD/LnNnVNwLob7s0GbtAefTEJfVJSGzT
3nc3NoAVtzP1Orfva8tD1v8wh5WQONNpT/4YcJJSQ2J2c7arD9D3H/DXed+FjM/0c06sFyAWquY1
sPEwpU4Z5sAsy3h5BIaNpvla/2OI0pnOcxYvmayembUilC5UxZFgCTJgFwsqNAluxMORFH/xZ7fZ
yJMiDydm+pDSrJ894WXQGT5/M1WbeoeXUecnBhXERklczP4WE+9FZ0lr+IiHGTkueHmQzL+8O/1K
HbyKmeHLaAoPRzlOxXE7iOgUAmzwoWUhHZI9QqZeKuzT6fn6FpUSu2poIuQE4EyGUGdHNDrYbA4C
YDkwgYxj4pltS0qEadmdUNxik5p+zXYfSLNeT7jzgaD999l0JjpiNt+V3M742d322D3e9oAKEoHL
4IXsR6TAgvUWhUqoZ0pzI6KIn09XAGFPxXsmQXk7i5rSxezolOuXbA4ztRr/ptpwGn91RU32pKal
IryO5zOGxkmOhzpmXxHQot6RaWxmRG1PuaFyNRQiGbuEFR6KPppyxdOaVx5eLGfdVr3BOUqoY60a
oKP+tNfFN1rZcPjpg63QdWe82/7HvJD+gW8AUWHI6W+yY/AB5SE8OCMhX3IZEq7Up4ENHWd8vpGT
uWGDR3oihRpH2W3nqC7gzOjKuv0IZf/uVYki+sEGhCjVm6gKdLQtxqh997neIbApvGClRnkDo9Bq
L1k7/O8WS2zjlAaiYrotYoVRrkxeMZVdnh2tIDR1elR2GOp+DZ7JglMI+EkNNyjR8ahMLeu/3goX
CbGlkTHlKq3p43H/8WH/ZObQhyY6tAhxQ8KM6di5Wj0gd95uXm3EqIQkpNaq/2g4dP4tWsvXF81A
53UGmX3swu6QHH8d45ZoZQwxUhTc4ol8wYE0S8yXJsJ2lAiWH4rEdQzK6Ox6eWcL2BMBXs96X15r
WcAnO2IRt7PoZDn5ZFLD7kmAcfsr2zgqaF/NDvNmq94tcLynGuhuLzs7552+4450Q8W6I05BHl5k
E8TIHF0I6BTb9nCWMn+xwsPzi57v5NA4DFORTYF/o2Rj/7KjGkBpfM949BbrphLevEZAgGUS9oSe
gb081cc70+LqWxRQfrYoTqh2aSLdUnpA06zAhmN/TYtewiq9ZEciog+Xk+7doPJ+te/h7iV3bDEl
lfqy1fK/ngrNN/Ccm/yl2K/MbnVX6z6sCXVjbsXhMq7kEDwrU6/ENmjk/6M/ZzBeI2xBgWtLyiMJ
m4dBPlagtrB1Jm34lNrgP9g5z8nxRJqSdlU5ga0kne1NP4kbv5rKAWow2ByBhWxXU1XVbd1+s+GH
B/AVu7JZfIO4JOT/1x9O/m7JNFM+oDgPBCTj0T1ImbQXJ+jRpb6kDLF7fS1Ro62Q97qMqKLr78mp
07Y3EXNh/UJSUuc22LvgRDCbqGS4i52QodbcE66y+sw4Hr03VOs8yMjAYZiME7R5FgeJ0Vha/+LS
QZuBKdHfg9x5D9bC1ZL4xvD46X5aOtdLH8p+HcB2D58teq7r5D8u0RyzriUCsbfZdVknRThQawy/
UeacX5+cQpNDgj+tKA93i2abGn8CwBQzqfldEqYzGs7FO7BzYKVU6VWKDozc7Deg8kmLirh2dN8v
BnlV6+0l1tP++SfJcL9pyEdG+Xl2c2bhwvJdJRelGmYt90UXHsy8lSZsbIkH7H7CY79f4UqB0HiP
RwGjoGaz0RmCVvpOblf5hAZYtluqflfoPpc7Dat06qx5avlj9spR0QrQDNltLb7Gh945owNYojzR
XPwf31fY589gpt0WDOMP0/HE4gmCeFqTp22BXa6cmqu5TP/WKw4uvAQD95s0cz9tnNIAHaozQIwE
FOWLbuu0kiqPsnbzekRdr7JbPVxjEbutEdn9V5M+c8iPU0suIXLm3jhV3kP6/atNdYdF9I62f6+Q
sdOsZ58WV06ZHMEE8j2YVj6DFp+mCHO0PVsQgL2WMNXX7g+RAtnHWegbkmuEU2Efxg3oG6ocSFD3
TYjQnTOdT4FzxGFiTzeUrzOvqDSZA8ZT1MvLAiipVlE1YcTHqcaJg81ZyBNqXbQaEdA5sJY3eciY
zrNwlVjBLXhcRVTCcRGl2W//mp+kzkQoaxSZ8DO6hB68yKSsbRV+ob6xm6KySTqx65d25b4+q9z/
gMaZxkJaNNkrbqW4gW8EwiSw1DcYKqRPC8pcXmR39uRHwOzNQ9+K95SQxwllcvC/QYeYtB3C7dT5
+I30aMbDxgPzfENNg1R9ijcibgZ6u+TsGFlG2M7YxlmjSngStwyQ2zlHNPRosQUyz5xxYkA18hBK
5TkZ7Zs/fqOdvtULAKqwVT3eFaSfiPaR0cWRKng8cDd6Uf4S8cta8c6dGUc9u6IEgtIVT8OfDEQT
j+qaZRYnEUjScTl3OH644wFkcDF0n6WdgXlBOF+cXJZq/RDcUUtw2Sv7feuQ2SZ3v2AWV5cMilbV
54KDW6DdHddFOS3DZVfPKf+mtbhAhBb6KkDPed4RSjUIjmUE8HdvKo/aNKdZaFZ5SrJs1CyFpS1x
AMjNjNArYvkM75jz6WXglt94UtGohEBpRvCmpVmRse6Kd0t8TCSmM+LbQcxzCwvdRSHJ9AU9Olv/
HIvRZv569yYzhw4hxnE69Yxt7fO91b5I1xtyJMxBxHsAsMu3NcGAdORvN/mLDWWA4txvLXa5fkCb
Mzs7Of/cu/VSQJESDToIzoIxL7ScOzk/ZrovRJVU0Lz4WY1hKGBmNz1JYrzvhSjcg2+ZDNRjM9AG
Kp2O8OsRrSX+9Wq6n5pubuzFx+ZTlgstgaNzYI3cR6MfMuh2ytLGk3RVV8xXmKn6lhKCGEsIcBoj
96K/Z+tyLmjUCXM6lWPnXTAiSB4bUUCo49rHWJvaa47c6qa8VeuzUdzkeIZhPY45+T1QTz0cbMlX
eWnad5SnU1SKEqBj0m0yUk4TgmWVxmOlWQ+aUSgKbt8+FJKdf8r/N6E1eGThL+In97xyfUb/dDfo
u4+XeSdr3oMoJvt7DvOE4N+XxL9BYT2pvZmRzxkEmvqQ9FlPYsEbs3XGQjER9Z/wh+m2idjU5tUc
TefZfAgCoD0ERLGsdheTNJsKi3rznXiCw5SGXG5CkPopX4e187bgoT2FE/YTqpxJg80b9Vx4g4UL
ayz9b1rfacczsuxXv2HyyC3IIiG2MCAJjKLiB/InYhy69Lyqi266eoElq4BSaOOMUCVayP5OeDxJ
LXQ0FNZ3nQePJoBF9a+nl1siVhL7aI4JVpFTghDnaOLfG4WxXPLP97bWJL3UucXEkeDf9fLxn2DM
5I9nJhS7SRyLoFQ8OH0ztpzRB3LvK6f5RoR8MmgZ1hwahGwO0bbvJzRGdjkjdq4PMj9DBrUouwed
STgD/7i3Qvik4trO2hjy33N7j1oXKoKlUl3m1VNR83bPnqlsTMJsSk2z/AhKVx1VCts8gJgSzyGZ
Jv5v4MU3+sadDBnQJXbyAYm/l6/eLKxrEg9nINX1aGGewgzYAvhEzBCgdWssdbSa5rrlV01mOQno
fHap5FZt/7GWBckSQ1T50CIz666A4+CXKW3N4s6NSoV4qqlaTge0VINqXNeoDBzK2YE8CzTmB3RX
4M6yy3ia9WsC7q9gwXqF6rlKlwRGOstEmWtVOLBC9d0eTYhHyheZWYhMgANJGvnSPnn7+3nT00mt
w0VUKdI6J1heKnUkQdE4xefSELCn9aa4jrKawQeIJO6k93Sa707dHBCa6XdkKA6rRg4xQrEFfogN
DdWWPSmWg73OirtBiyTs2uZwpR1CW1+1sG1DGP7YgTak/ERDQXBVN020ADzNc+WoT6bI4gWCzNcl
zZo8LVkQGkEdZvOpKB2a4MBPvNeEw8Vg8QzIYfRDISqZ2hRk1Mo7BuLEVsk7iYSWs6AiaZBGwdkG
MZFUc01ULOwusULfaR1BzsFy+kEKudWZgpTIWZ+W8AIVkfbrfQUpUpdVFrsGRgUPThnUR+Hp4hKG
FHx0N0WSplGrPBcxZiUO7R0dFP4J5KTKFHqcBCwsBip/hR3p4K1AdgFYmFFaartp17I5FXdhdeIA
VOlDj6BBDOdqnGElICt6wOdJ5cp5sgq8sMM7hvIahytpWgfVt1oc7IRTv0hZtFU3lZvBgKVnr+m6
wVxHb1QUyVaIPCfOp6DowGt4gOmgNK1AL4pS2N1WsBG1WOOWBBUZ96XZQj5OXfaOS9o7R/EPVyXT
i25WnHtHC4R7kc/irreC66qpvCcVa5gy01z3kOz1LCZElS3/Vs5vFF/uxVO+BhD76iOkR7zM42d0
jpjHGrcC+WzcclthwOfzxjpADH9tUN8H7JmxDtUPkGlRAMKBakQcOOINU7b6A5jnYviLfJUWP0Ww
TbMVvRR4Wf2OdpRtrM4CgY6gWMnRa2gBXyivr0wzs3Y2lAlBChlJ9jI4Muk/gc0p3QNxRyvOonm2
mlDK75/5bIoggAALOzJMzf/6DLbNJmbo+EMQVL/BtDRmVRrWtppavX9E0O/Uv3DO9CpO05ftPqF0
5Nts0qcMdL/h8xWKOLQHhU2KdLfMlATkImQQDdrGDi11F2+2+OsYFkcCx+SkO6cb2Hbrv1yaLUiI
hcZ47lHFFvHr89T+krEchs/c+zdMY/aP8MOKy93+l+vMz8RWrbqy4PcTKYZYEgVG4q8CRI5/RssI
HLIaE6YbqzAjmdxrCohZZ8u8fxZKvbUDpmmjfNB1Jx+HEEhx8o7rZft1IvOTOMvcFdKQa53iW1d2
qBEEpSTmH0royPSY5NHlmzaCNE5xOxYFJBl6Tcsa+07m4H0mJevkjj6Mv3MJ4vN4O6u+z10Skiiu
p2q4neUGiRxRIsJUvvpPb8b6SWQooS1ojwIPYvMozFnmvCGpcdtKpI+2DWmrXnzv+uSRDQQIkujB
uZx+g5QGZ5Bgq/1Vh1HzuQWexDO6KuayrljK4iHCWUFTa6xi1PJyXWvQdd2+9P5rp4e8YsGCud00
Z/b7p8Jk7c/4Gy1HlpxcDsnLykcCT+3/+Cb3Q1QN95H1vjjjgeSRdtBj4hUvJWMaCNzZXcFgxarH
hnn0d4sBJHpTUahecSOiGFwWpfDEPzjZS/RM4lZn4wM3F3ptbhxEfvFIj++YdpkERQYggkt48pga
m3/eXQbJQmx6ipog3R9+ATrR6qV3WVti32UarRFca+OKg7NiHeId+7A7kKWWtvYMjwBBjwBWlTzI
2LIVNAzfG6JcTMTH+gvNuRh8bCkuqBEjuj+ZxS28xqOt1DcHEFcLtY6xOaYEchdmwcwRkLhZjQ6k
Axr5fwMiiLzZK96TRKlBGcdEKWa5+KUF2hUFDJMyxwRnEvNPABbJZtorLPvk+LroLVVswido6QHm
jb8IsBeHIAV2i0qAZp+hxbMHt4SXgsWn02bHUp66/GZ0RN5hznUm+C9sPaDuMiUXgtQR13XTYhSI
QN1W2IqU9LsZ+2+zyyGeS70y2eD8+gH0hWVHwRnJvbET0IOrEdUhC0U3UveiPRlImDp1ChZ+NIQN
lCb4vorqqf3Y1SAT0P5C+MgwBNZRcx8SocheVafTYSz+HZPbyN9NEHUVnqD5i9iw3ZjdQLAv1TQa
C9aSKmjhVA1YNXZPRkHHHPfDxnUgzUkd1V4gvBdBDa5ijDECGCRZDWcfqQG7m5eqcfZw7FTOkDaW
S3ot7mGYUO8N5qCZLoI4dstDRv9AdIwdRMo7OhWDL82csjNogz4txsuzpfb5V8Muj0AAPSkIlXbT
7FF1ngnqf8rUk+D0DY45quusAKQPs8vKd2xRJTKbLlUKGcSW0z+YaXV7NE4CMvoYhJYnTTfX+SLe
1G/jMuzrq+LMBJfqfb9RgL925lJBJz8E1oZHuupS+gHkxUqgcyasqSeXL7j8nm7zDGkaMZPnJHDD
8LJoPm9cecbTPrzgLQlo+mLw5YV+3p3C+FoZPNbWWwaVNlp04sexqcNTP/PT0pBKMmEbB8igEgEd
+HAa3GaMGE04GeXmKu8fCGHiSgHLsdj5rZXZI5IC5q9dWWD63d8XZZYyQ7nN2bQCJ4B2qwmHlzCp
V37jkD8OTkUAvUrTftqknR1r1Zhv3SXR4Tdo2usLOwoxCAX8AMHO7nPruE8hfADba0AGVA2Fb3lO
li+iIPYuSHw0xwqFzwi6yv225Hz18HB6c7VeBIvRQ86ON+WzDB3Wdt/x7antI/EROT9LHmd3pCzV
MBQVhLKaXZsd5mkYsWOA1+ouU1WUyh/cQ8F4Pc/ziZNze299adqhFPJoSYlalUDS5tTlVUq6Jqvp
RxDJciTAIZtdcwAVI2E4sYz7jP/TFJ1czWHmVmG82Ka2kpBK39qTOnge/eQlMGyq6nmP5I6utgaJ
LVJb8STI3UIoiKfHz2Y9IpSzU084CRQYuED15RVB3j2lo+pLXxbAhiC3cnpNcQHPISbAvmLWgX4S
0+le+BK+Mil2EwOLbOPqxvvm+k9+BXRxZsopYlTAFKEOZd+rKFpS69Pl5FfLYW8MA5Ihlxc8Ycdu
NKTG4SC6xT0Mkbmae35fqYeDDvYU728I7AZvAqftyg6mlgnpoQlSf+cLpWcPmRsmuuULaI2WnGm2
IV8G1WN49+zFU0Ct5uJa9wzcyiBj6xw07HdWQVodqZKDGcgEZKew8kekpNWpndMZuQXngkDg2Uq4
3rY2iuI0YdpO5IxjKKD3phFRMJpe16ln8AIrIZbxybYgSLfOAG0chf36gjRcMKQDZ8sL9Q8jVv+h
WLAS1ZWRgcfEdvezhyNn+1Nz30CH6yxf14HMmp5uFHDRTjKJHjsFYHNWEkSXsTMIgtdSNz07Qqo0
MGZdbO2/5Qq4QYHdD1MmKgnQvoI09neltg4GiktLEyE/7NUrDGVbppx4tfeuSQ7xEaiqlGfotvDB
nCOYLe3JLJWd13RbvDTEI3RknDgbGvdwQ+RZ4//bDAwZTle5VVUdLLMNdiB9LyHbtNwfaJGgTPs8
YnJ3ANZ8GAkgxwkI5SEYQ/fUzIO37A5JvEhfDiOALaVR6BMmv/d6HrKJBEIjcIQ/ECGPwUM5emPR
S2JxASMYakQiW0LKrLvzktjHosrO2DggDD2oBK3CyBTPUPxS9YiV22Dcd5KkH0jaB1DKrFlXEG1h
pAkRvmqHjkdXwEJmig1+Bvx0Xe9l4cB9HBu2J9AnvcJWji7X7DZM8ow4JKz//8ZQ8FDNmguBaHq+
7tooRjGEhZFsFm1iwD4Nx1fp4+75eDBhbfduJVjYnuz6c1sNyTI71pkppK10TRtrhlzeokkDWV8f
f6RJIUUBhYXJAP8KRmentW7XynHPDZQ2TOJkEql1sTsVv3sFT8KUCgYuPX+3OWu3iL04a3Xq+M/t
qJjjh1lI1LYVsf7KQw7ciZtKHrzIWJDUKR8Iz+Ra7bJIxF0K8vRL41+vsPIEiUvcBjrTWYvOYsAc
bbpl00OwgIhphmbj59uNTVVq+ZYpytp8Nf6NEk6PR5VdcJVPAinrkB4acOOlvFOpg2f5T92Avyk8
LoD4D1gQtWhsasCHBb1oQAXSBM/n7hwlVfiYl8fNF4VclrM8/Q1br2b1OsuXZa7xrpBW0KU8XjKW
nP33R5nqocXK5LT3cup5qBXOvKQOcl85UX/Sfq0jzOEzADUIhnjFkdYM4vPF4T/ITn5HHvvpIg1M
uqCrgVSYh4mxrr2wAEAv/MR7z0PCyTIkH42zSRHa1uEBRhTAsw6scHbz3cDq8QODf4BtPYZWcKCZ
HhyfkunYjyacULOL8ZDm3xb86qLV5/L2N3BFnCoE2FwgfsDx4+L9+uABc+/IZPzq6AUnyJ5fRWq6
M06c/owhHhUxeIp76X3Wvgx4PrUcgiCZOsvA2Bg0ha97dPz4e/xY9r7kFml1bQ818DsdeLPjmKDh
IGn2CryJfpc3lpMz13rjfvGIAYbE/jcxx4xBVzogNoR8LRSUl9wbzr0Xv5U1iViD3LUH0HnNnkdA
8fDc+Vi/01Xbvq3lwubZx3RadTFUs69gG5Zj1uoDo/prdfMfJm16f2kZ2okxWn/TU89TAdgeymIu
FMQYqI2RvTM/vHmTd1DKjHDDTqFVEze9yP9IGWdm3Nd4tqEM/D+LHGEMTU57lc7MT9ek1IwgEXzi
v1TeIRvWX+wpjRaaQf9bT4lR6b4eu5XI6/c4yOctV6cPJsmr6TbMK6+xOzLVlo6tlsvNi1/mKx5c
oiW9niqa3ANhQfAzqQAv2izc7rFRAms85LGGW6VsdFqudQH6+ZjJpV+aGNReX6R+pl/scPcl6rET
Me1Po8JizpXDO53QEKTByRWITlNMGJfgagGOQ0bNxW34GFCfvc4mlqNFYT1c9w9SzncA9V4K5Yo1
eKJbfyRpC6YNFNvd4JDbgTVM2e9c5nJHmov7a3PV0eMTItIDy0xzwybUajrGreoam/CK2PLTHEvr
z4ew6T2HDozMie589HSEoXePjDTJ/wNrL7mK5OQ8kltusByy7ttwCnSAa0AN5q3Z4F7zjw+kfNMP
ivKA8pLC9Hk+aSiFaTz88jUFGfvhqJBOxKRoR5IX8JaAIP7OKXPfoHSsj7gkN/1R7m5rgJdEL+GM
Swwt9XeE1iihg4vUr6thoCX0+xisYkTZ8fr49XpSJWCfCkbyLXN8snUVGTjbBrcHWTNXVz33V0/J
QzObuaw/GIsj79uSi0iTsfR1ytkoSqsj/bdTCxrN3aSdwoF4WY/VDVd2cFe6XkQuBlbYLH7hQtre
oNSClH9eotC3301rxXcZS03a3MJ94YRPUzhqD+JbGh83tUiyNe6+T7wuz1eW8Ol1YEJVVyAlHky/
WRN4Ue0/dzeZTBeLbUkL5hXDn0DtExBph8c3FlKU2dfjIrzrJH/e+FvjluJTS8JR89pud7Hn6uNz
nqDwKuQ/Q+btxTZVlhaT9sybsZf6XjOU/XoZLv91kfxzFo4ie8eloQHLEPfqpRe2FU9kwxTHmO9p
HP6o9IMufTLKNZSrNCe7w/AV0YSLc6I0KNdweN8T1ENslSY61/OvXg9oGgZCDHyA+kGHlGdMvR4p
ypKCcAtJqjD212jd7ngRjJev6gMtLSnk9St253CRY21GJLkzyNvPOVPAbM8JXEDkp967wYi0C9K5
HeBhlYM45c3YhA+/PuoKzkMM+r+wtbdWCu53IVzrnyDdjVMmKPlaYuddCwxx2/1rSVqTi+87iIMI
XjFV6WTv73H9Ewgdrd364C00OiZ1XAfCH0dgztrYUSwO0MBx7AfqzFIW0BHK0d+9gSZ7K94IpgfA
5enS76Jl5jbW1/QoInebAftYjrUk3DZS59KiPNrYb0gMgj44Fo162ZWtxErsE8SIYm43NhBQ6JHQ
mxTDS7Ncbo2FDOytXYqyDhiWkIc+p8xuqFW7IAGVr+kXPjHOUYz3yRPtP5vDkKfmcYgDnMVtRLRy
2D5OZ6knA06YBEHhTnU5fEyLUW7G6hMHEgdWGuRbDnTjoyet1HoRZGEQDHrn5x4V/oYRidx9DyO0
y4NSrjiHsyf4lp8B73hPP6o/aRDu3uY/x06R/b0eppppdK2Z6ltirKJObLj6ekWztCBf6ORG4Oyk
3ZwbWLdGtWKcOowRMkYhzblAK4O7oILv8xGB5Af36RKlRkXKQxs6+oVQGAhwGXo8Tq8K0H7poVTI
hybb+n6llM+nlkEn2jB4vgIUIGBjiFg1V0CnCnEaz/bNS6CF1xTYQgZC3X9PvdEfjAWlNe7Uw9UE
xXeZbck4tPMr7Jkm6He6Tw/napzW1ZPX+DH7h8YLMSvnUOS8Mi+87NfLqJ7mLjbuGKthp8FILnVR
nAN3O5wdIKlczPb2QeHIoBh+bGv071VzRPi/++fucN2MZ9JjxS6huL1R9iOswA0bYoeghkt1CZ0b
RCaeFOv1MRlXTStXE0HaqajAWzn6lByQdmPQAqSXO3fx3q9x+rmodUXtrIwJUq+0eQ/kU2jkw3Wc
siKTdIHNUnhFgngvimBNMGBJIAyLj+Pa5k4rSyxqNInxkX0VhfeHIA5mQuooulzcnPP81M3j1kT+
vkCmnQlnTf/yixEtTVRwMXrX4CNIzyLgYqyDWOBRHhxiohFxyfHmGLEd4cYzla669HsBgLWvwH6a
baUE8fO0elLoXk7Pf/sMa3ChQV+YDBZa/kgmptJDzjNRmn5i1OG454753iulVIUUDoW8EVhKZMjq
Ir1QlRoVpaOgcBL940gRHVo8lG4+PYzmR4Juic0uMMSkNjxU3f2huaRNb5vXWSdQmL4fd3v+1tdj
+CPh3t+Ni8FKxnSB0IXuGbdW15E+wbtUE22l2RnCX3ZiUA6RHhYfZrmxIPS/YI/UOhBSvJrRs9n7
v1IHFooyw5OfWua3Mh1tlXOxG2AXukpN9b745svqNRupUVMNXrApUAERHhx71Rt2wFrGWai+cMnC
ClfbWw3YRt9AJPimq+y+hHprbNu1mN6eJs23EEqenxK1VVgPpiaWbUxHpZ0oxW/mDiMF3IgIJXfy
cJUCbCZMjH2jJY2GTeqV8SkmJzBptKFCA9/fTv5RCrp4OWjc734DIZig6zOb/2w6a82VBkz2hRy0
c69JXHx/3VTHq55+3oPvxjdx99CzOxSQbdAMlATZbflcEExdGpDTI0W0rIHtU15GEiKxbm/HRnhl
3GoBf/QSKbOQWD9Wn8XlE+tdoAJWv7imvKgdVT2289HPumGlmd0GXzpLpbgUfxdMN+HsffI1EPIe
RE4RaYlVmwe8ozlvbVhPgW+XTGmXz2MirpeW4gO5RNAfHQ5Aat5ZqpGBwbyaDzFA+eTe8FZMXYXe
Ffz6fKSKUUbH4qUQvChGsVjVq0qrIWRNF1eejdKXnY18EM+EdqcfTAnMq+oDukZFvwnBuYlH6M1v
5xHLrzDJDTsQtap2HU0ToVrgcXg1fdjc3eu6jn79kUnVE/c7gP9p+jbdgtEq5gZ0APGh3+OICrPY
9Iqc9nTdIz+gdawe2m7zJAcx/VrqCaJleXyBHWOqZxM0pn0JH5mjFo1q8b11fodqdOvo/hOn2ZNd
kFj3UuFJ6+/3LqeJdCeFydNra7Tqlu/QHjqWbOusHovKP0q+E4byoFnfVWxz2Dp7h/+Caod98Yqv
2yYVdNd4vluUlt5sIdjgqMJRvS2x+X2N8PGpP7PxRoragKgSGrDYVWn2o0YdBW2AmrjabWUWH6VO
yWADMpjhPmPkxrdTA5NxsPlHyTlU8z7y8HFKPyPEteO9nh+0wSQ3Y+hy3NYp6Htbm89g+loLWzyl
qhdBAQLcDzbCGzlWYwgjS22nlkGOMIF7XFgM70aZ8Q3e/soLyUmik8jy2pfvQ7EupBGl11MXq8f8
oDccurSaMNjbL8K+f8sNgcwWhTFIBcFKDf1rVe9HMloVGHWffPC2NKz0jL4L2ozUk6yDMwa6cQPb
a///8CAbZn67y0F4XKPxR53wWihPOX6vAO8pazKnMsqSEkspP99zy4KExb7ijYXIdLJ6aFkU5vfU
0OIeTONTh0zZWrY9PcebLepiDahmlJ+BdqLe3Uljd3T0nuqUUJt/YmtWxfzCsbQ5a2/76gBo2BC3
rCNQC3pCBdRKBY5tuLM/+Dhs2kFSAWDSqLjKq+IrY7ZBIZ0eV4h19R2fhYx2ZwzmXcZXPwiEqhi3
EgeXkp3c3U9pcvY6NgYsuejFmTKjoGHpXlKHid5R4Q44P/yoT0x2/zGGv5utX5rpW3vK5DMwKo4/
OndteMwKY2OUjxposFCOc39HxtxvJP0ahu9vrzSamy0P1ihCMXoFYH6etlOBnepWfxq7s/CI0Rwk
bhVcGFb4vPIYFrHgKqjj9BqMivLPpryrI6m0S8IcDfC9/d710yO1iHenekC3nA7b1IWR+Yr85ruO
Dlakpl8rr98iusgBGdlo/DBCmhTDzgXAqzpf5UhYH/CjKkdT1pwl6CnCc5qwizSIVNbGIfm2vdCm
Bf0NT5Xyj8xXQxByXTmZ/hn1UARW0eWW6fPjCPoONiXRIJvFytB9JgSYtnsmtHE+UL0ev3tlov8i
H0VGa09lvPmDxS9Fl4DzcISSz28zmQrsngEuhaC8jc9TDD8nKxwwMSwiGOuJ4/45F+R9hsUpzKaH
DMCcnvsx2ampH3AsoWXgta7i37Mu7FubTJ/i5YLd1o+F2pnejzlkkfoow6uawHcORswDVoyite3y
wP1QYACwbRNsG3eJWrLrOod16CDgeJjFIQHh2v+twf1d1m/8mC7lIt6w2Kffg+di1c5O1/n7cqN7
KuDH+gX8+An/Pn5nfIN7HSkegCXB0k72RTytiL6xIsW1VBeDkdQBGLE48v/TMRddf7gv8JyV0cac
Lf9GEcCbvDjwuw5Co+7HEjALsY/+0d5U9dreuVAVyhSxSVHRuAlZTu4XH9kKwKcTX3oQFtc+7K+V
1UNq1ngeDkYpSj3T5QpTX9pW45mAeehBE47qCnxYiN4UjFD4kIqBaBwoun/pKKeI/tlOMwm/vvnZ
9Z4LMJlCK/c52H6QYy8ME2vvQVZRW+1+XdVJajqT7BkXiC5s02KaTM4jVnKnPb/jpa2Y2hzqC43R
JMRRY9lYFig/GnnbGrpRjkqG+UmgmLoVat4HzUHJ7R+AMQjktyyBIcmxRguk4b4px9L+7Je+WlTp
s3zX/yykuACK1M1p+vbkjKvRcVbSyNiReIxwxBEqnVk2sDSZU3LH/ie+Jyk5neX8BUfTXlTjXEX6
yulrKEpdos2y5YbccrgsFWUZ+yMnvWf/pcH4otzaWnYDZUAnsO0UXPgkhTagn6tFJSPg5iYHT1bw
JOg1g+5LdjHJyDpecyS9vYRpT6aKo6/VFVjk87yNXtQnWcV5QUGCy98P3R5GWg1Env9KyD2f9dnM
Jb/PUVFQoZ41chJUTyF8s+iTwD/s9OKl25H1u2dTI9TQT5zrnc/D/VEY17yA3mf3C4RumbuYcoeQ
rJxAguVhQZc1SCDsAmTUgwKKEynbPeKtUNOHoxFU1bIEQjYPv8Z7IMaiXj0bvek256Umd4Rizh5h
IhpVFm7Q7CoUK/H1KhT7H9AeZX11Yb3V9tueRFWdmaLupJOydUTMx7d/Ko/4nNGYaOEACTgY6AGF
t6mDVB8Y3HkC+SCP68JS6HlgYvKQNYPYac6EuWgfp9O5DWE76Mhk2A31hdVbG/HWVQGj1yzKE1Ky
wBLStor58mcPFD0YSzMAAX1hFsrGUDrxrZin8iMWNN09WX97ksSrNSjO3si9o67MO9NYn4XGUU92
5lXZUCv696YDMfbO3Qy54XO9l/wMI/clwrDnUFhTVKqkJl425Dv42/g4gZyVTOemeNfdLa6d6zoG
MTmZS0w5qyo6KLQ6bd4EgI73iByY8k51YhAqFgQc3Dnq+LSg520nenZrd72W5gZ8rRlfGkCbI8UF
KgtkUJNnl2uO76qUz1fSrY0v6zsrmt1kUDp+pvm35RTokROGMvCtA7/TMteIrJdGec16qt2rKzSg
S8cS5uRMZTN6FJqI6lGkPlExxLkUShNmXIfWae0slZ6JJJunmuiBG+JrX1Ng6Rmcq5xEAkOieqzb
XTGc6yxK8w840vgvguim6/iFDP8fYJ47RSPMzCMag4xLu+pSWN5zomKZmTz9njYiMP7OZbia5cqf
9LhTYA4bud/qYqshEz5X78tRsHfim3E2RIoZQ3opoUhiEj7AmyWZD/Edua4Nu0EVd/SrUDMgSe9B
wEIMM3gaPs6ex9ic9l5nWKWqBdeUvwkE7dNDqbxZhvj4Qaao/Hk4L+RNqwfTn8IQfSf+XstwCbyO
yGOfDSVe1+AbUof+RfXYzrN/Kt1b0GxO0wXHRu39fVexh5DK0Ru6J2miRJ+on4Yhu5qRzx0A7sua
GXIPKRxFoexg3nTbGZoGkaMksWQ4+JfEiowS2MjkZu9ev0CyOBDDNsqJuzsBEPrOjXEgHZn7VI6d
2nMWkMZDuQ9YoyTERAby63LllxxaXumb+8YOGXcF+/wXeOihJc2gHdo2qK7/1ApBt6x3X2SiyBXs
uU0yBfYPva/0NDTDkR7p/bNDkkEM0wPj5uAAmKsZ2s0jjZ9/ebNTSUHdqhTHo5Df8MDlJtqRMF1/
3xf5ouBvukbFI7ApBsXr2+jMwY4ODDLqYbbROjS8lBxvkTGf0ZKs0DynJUmfewXguevWqOpY6N7g
uOZfR+YKGpYRSXcJNiKJkvkma3a3zB5YvRGx0zDoyAGs4s5ZPl8iIh6Y5nnPIpdLSUKPZAeHa7Hg
OZojLICVlz9+0ZfsWp3YCcBkU+u5FeSmVoJ4ilfiF2nsA7SyJPvvnZMVGv3bjkawaYkkt4e6gf2t
mk327u190N7/lIp1d/tP+Lk+t0vof2W25r+6A2jwY1BCelYdcV70tfoB8mzS+QNLeko2R4+8/iu5
qzSTNnTiqtoQm6XIrvJ4yJBi1boPxn6egYe96JmrgDAvM3hsyTfM6wx1209Csf+LMSrJIk3/lC7z
SgewgkdVHSOZpNKJHKYrhyVE8KeJq0h41Qhasex0G0SsRbCwEuGpoo0NaGZFObJS9H/Nys18jT0K
y9WRRAFZFyUbDziby2m8gjzl5Ni+/zC9wXpJ0tAjKDbo58fr8luhmw00QsWWprj3JYxeYMk0xCC+
UcaCCwogJqwSRjzWM2K2Hxc5z091xS8zxeIJX/IQcwLlQdm87EzweKRolupWip6MgInaZCj2yzms
qu4bGHZYYGIlt00BOBnpiCnuTY1b+jzgHd1BXycYapDFduqkqh5mcJ33H/FpSESv+NDKx8NFJs0v
r556VasJRESZvrM35qLgHVStOhrbxAM1H+H7j5yZ0iKT/qSlHwvPV5M0JITBhU8DMYC0KIOiFkVz
WmDDHJ18uY8BhSHgrHf3/uk4WbsLsoEw2JAJjAooOqy+6DNKqo/AP5mTkS+7dcRnOCEgKse7VOU3
2LZAFJL27rw2gysd6oyiunYGxssa4fcEfHf1epWnVLv6MKU2J0iaw7/TdWnmlo+rAtIF2dwFHD9y
xROcMhFa2FP54/shvJvBonhGknsJT77WQtdW8fzCWQk21wNilYso4oe+GEUUbwNE5r3t4SMDohh7
E764aDGQ0nF+IgCVP6L0Z+DISuWP62qiLxQ9A/N3oo8KpN2Ipca2SL8y5MWmrBbqsDazKSfR9nLU
ux4OAhC33Ln/25u+sCAYwjmDPfU6fqfHSrpb7tfvTzIzFDsKwCzPw9Jfk7jCvoaZVBxLEV7enPpk
/wb6IRG9G8UFKaZ29ElzFBwIw7vTKe0AO14cC1LrJCnmAoMtHl8jzXRPziH7MFzFDk1rqVCSrrok
HI5qaJYeMuBPv6f/MuIiXUS+NpQrJ9ZHJ1LlrRqq+8zTlxmf9zgpeqybatOt9HZTokHlGNWYRCQU
BVmbrADneKDBCpXE8L83SEflEOdUS+K7p/FFuZKfAlQibpb+gkVcfUmkYR94bvc5ch2r0W5RH5NY
5FFIcBacLN4r0H2iiOOxxN+5v08XEVaqYr3uxNkra9zIqEI75Zqf7gmK47CULgq6+5COryugtqk7
pDgmlOK+ER0hJ5MYYyT5+hvCnd/TWDMWo4+m42OEUIM3rsIivPdxWSKFGUup/HWG6tLxiJzELbfU
a5bhEyKN6lOBZrD2KxtM0gsGrwDvsRWDQEwekkfkExKko44xrQ0a5vnWQa6TkEIFZkq42YPp32cF
xjxfmUV8aqt/SSKSjJyWWqzIJ2BToyzCktBNMM+wVryJnMdojML1/ZSP/NZvSJawUJbcorRpSDV5
eSRB0V/aNXO6vwCqMrbhU+RpfTFUgmpXdDlY+7lmyQdotxvO5NWG8BXLx0CDMaTcTYgp8pE/eq7y
hkPJCZp17XIZK+aDD/K/NxdmybivlU8weh3koA4VpUCHEKAo4v6EtKTYlASOtyGDZG6Vrkjo9Mml
AGOGV2qiKh/b0szb+8MHiMY55EeG2x0xHbooQQwrMTYCdxy0ZAi7yS78f0vROvQcOIQQoFg7zm3Q
sN3ORSqJcbtYesMCshEShAKtwIk9t+9UD0kADioeNifonW9Nj5pdEzEwbdOhd9i5n0f0k0EhQ4Lz
hw/O0Aktv0aFa2xf0TufIaNCbeJXKegt3KHgvXrTGeFngJalxX2y24x40tZmMnAKgFUZWkyM0n2r
AWAz4pLSi0H9C8R3wvEhPvjbWM1SDtdw8M8i31lD6NNPeXK31jeRwbtmDhM09g4XKo3+xuGYBG6X
CVocnEkNYQLPqWt1KtN1QRxjI7iwLX1eY79ky3wLtDfgz5tC28J5eVDngNe7n6lUYBX4oleo4hyy
S2+Oaaez8EqCy4ZcAeyVy4jRdWBrp+HzA/yeIbVbnToOfQnrZKrJ315LuMLoKtF2QFGM53sH/EG3
Ro+GqOHbYrmC9Eveb4Neg/eNdsRgcpLOSJ33Nh8hmTAueHpwsOx7B1qLddRqN/LA8Pv1Wc7MwzZd
B83LtQ4AcEzSG/LJBBgYHl00PEO7yGuAnWZdiKzKMXZ3ymYO0PId+1WatZn7IPnU0PmrEai7pYdw
ujgyB3F0YoT9w35H2ZJHBPtANz1vNDVI1dJuWtK3UqRwwTN4MS4DaI2t2+4PfxPwPLKSYDIiNady
zzzW2lOrNLVI+963bhunbbbo1/hYSTdmdOVxCvkE26UcrNiIGcHAhHL88PzrPbckOJ9xuHnooAUi
I6bx0pEYJocPTBpst5WKC1MV+FeaO9ljSytLOws71dRIjQKBe/nW2O2dKeO5cLpPKiKUkadjLhuN
/cr6UUNW5mV9QV43xmlUMpSdYgmAdNgo4KBsfCs+aDCrFQLTFpDXZbqrBNF8Wxi6JHrARqmu57YK
JLoHrzgx50shKcGenxvkA8YaTaZLRBMpfuWnaVdYLiC1ftN9BEs3JGvzhWZJEOKBiMwER+CyhvCl
ojYiV35UYfq8x8wxCTw0sE46wWM2jRpzxWiQ7RMogPpzDq1QiCfjduNk6WNHpBX0pTEZN3bz2DlU
zq36y2AphS6ikDyiZbiOx1fMGdgyUqx3G4ERQ07iN1u+mHfbahItq+RNo1Gc2sIuD1cyErt4n5jU
dP8oEeYRnbbEjNsqrVL9jtzOS1qZ61miDApsr66+V1mp411agSPuRSQ3ZByOuTh+K/MHCeMa+Rof
0ebiamzP/nJcZ5GuCnzD5BhInrIX/YKMKvHt/n4J+wnL7wWqWEieIR8B++hqj8lmWb/mHmkvrqg+
H46MpRWoQsQ4Ngi7YucNDjVHZXoLv8EiDCY4PNT/5vQRbSOHWXWf9IcAJRjhwKeBXBqo21oDArjR
ke85HGW1JhqinkwgPagv24772Btf6ROBBQwFiz/GvE3M/vQPvKAuNT5JhzbzyfntDB8C3MpRO30w
Z2k1ySkfR1XL4SRG/AXF6afb0oq0PPRvf2p7nmuXDdhr45fbo4RCn02f96C31cmKFzMhK3/xTKz9
w60qLVLMU+2YYyoAO7y7mDb/oAkppdfEwu6TY3gkVlIkIk0uuZtHOe3e27OoNTs2fjl283t37zKa
DVqd+FiP80h8coGOhkMCZ7bKx8h2fTOfKaVFtyqUCeb8hdVryhOOLmpod0sN2E+Lhl8PnHNjDmKc
n3izwa5DI0CbDzRhzPUBb5vpa/tU+fjIzI94aO2uoabB+l0kMa4bxY7I2vLLoBXHAhh9uERfAMCQ
nVxfo5UlbDfZSoQL8j2OwnkuDk6vx9slMoUs+/thOB6lgPbNTdTEQfx1sRMlU90GT0TSrt6T4HQD
nz1ZdsmupPc46u61VskhRBKGrITeHFc31ywSMuYFjlsOZ7iNqHFs1y354yilJbjsBUNButWrqCAZ
Wwd1X7RrM9YrH4hLleBDxyEPx7StwGfJMrulpTT1h1O1FRx7PdXYzZPjYy6F/IUcKH53VOmNFJ+4
Fn8M7atmBJng3C3rfHI8ghjLD0p/TvHGjC4T3GGDHiFT9rir7XQXRqFtHvg9A+SfP8mYRbf0sRM+
6QsN5NM/mojsm3Cxti1eOd1fCbP/hQKpDNyOqTDlwJJ/XpEl4HmqYI5U1EJleSo/B4qBrBqY9l+x
1CT9PYirmpEgIczMYhrzluLoMx2CDZdWE+DIaq9MfSa6HSSo935WV9+5W+2UCyEd1d9zH7o8sXv4
ONoKke0eFGp9hCtwpIFxFY8n+lJ8DfFQ2iUSkqzaPZCQBLofkyLt6IW4Qrw4OqdPnskZf00xdPtB
fGmI5gEb5K4MALP1Fh3xzmHeTixWzwoiv+Efu9csbmsY7Hssx8QvHLWHx4OxtNWNwm+paS7kO4T2
KAqKRw3sHM0urFgmkSt6P1cw8gHwDnJ4zoQyEL/gXC+YTNoSOOvjBAYarY7mT9OXcA5YK7RxL61o
csk5jSCMG7UdGJ0WUqHSxcqMUJTGgSgKRa7dVRY25Q30M0rwZKxmayGOIHpKyiQvrmEEyyigsZYq
wtff/ElRMMgb9ppxXhcAmApL0dbqKjHa5M4+74b1Ypk6ZZyvIcu1vw1UyEluPxyfsKrNwq+m+cyH
eYg3yaH/V5upojSsDppoKSUmuwhiJAdKr4DKQN6EHMJSxhKy3xgsZ2Yi3Zt35Ux4MTR6u0wN5Evo
diDiinWmoUpq0rG9l/wBLx2tXaKsL7nMLY3cgxh8Kh0qBhgsoQDX7WtsybqsGlTIDSpPoM/rVtbS
5hjQOPwwi84C+Hu9AUC/eEgv5wYxWxV0JJS66vWy5AiBAbsFf0qpH64PJ6xOvnQKVSS4a7Xv/ddx
zRXCt4K/lHRbTlZK1Tb9fK9EaYV/E5j5nSNiqsrhBd5i8zmzEDD+3fymKykiAm2a15rRSyMsK5nE
am9yK971XVa0nFcoZgaNS9Wbg54GFt54SSnsZyXeowfxuApqTCk6QlU+oDJ2yrU+k/lG0x7JgW6L
6nlWx8Fm8a8kz94MMwYEffVxab7bBB/2nwSCAgDiFvHZVSy6R7eXowZ6KqNFUJ7UQYx1WsYo+E2h
u8//rI1nCNCHPagBLfdaqf3NrdqPGmD/VYSJvhGEmOms/jvSbN7XbQR4j4EYGafGVh0ApUwV2qKY
PF2DaTayI72slqZN3vw4/MkBd/rVhWU95a12MkCw2ChDB+EcDYuF2iGrEIUajdPDDiKrEMuiuN0O
DltCT6eqooYhFPfo/am00mo9jDgKr3CCJQUtVdyoBwtVlRu/ENXahzsHjEisooWV2PeDo4iYlOcb
eX+s3qNbJZQrXZ2pt+hX8nBoe8xFJDcORDSFIiYJq4NikcsrFpQkg2BT8q79KOWOQA1gIOnIDs4g
njKRJMkD/2J0Yqec7yTSKpN0eQ2T0It2XQgL9XuI8pn1HuCutFlIK6i1JQkZFjrgOzCUajipU8W3
x4ZC4GePlxTT2TFApxsQ3LgWwB6HySYZLxkQEhTkqTy91bSZfkL3tXYB7h47RboCmzRVG+jD2pkO
k6354Now4BLbNK13K/qAek0YMA1o+A6OJPNKf0PtpMNFLpLJJsnOON2Fyl9WCypHeEOCPy5ZONmH
U4/YAWUT5YvRd7tiVUmCZZnhD0OI66su8nwFi3vWoIaARvSaO8F9aTO3pKtcZN4B430E+tYklgOJ
k0F6bZ7HZS1Q8igW1IV+q2oETnOwG2FcCSeNctZDN57YhDE30BbY+quIcbcsTJ6QG0YffnE08y+T
KLHUv8DSf5GmISHysVZ333mb/qSsSvhtZA6saoZ91R2GOIIRyA6c4BUGYwRlA5lgEdqZp3+8CL0L
MzOostY6XP3VobVonOtCgEOYAsg1quodj4OyWYEkToolDbtcaAqWj1lOx+nSNY684Y85Q9Ft0vO1
3Z+Ih9oTCGrH5WPgWP+ptm6gZrYlylTCzRD7N1a88qwXi/9GPMmXf2qky0QLTSl/TjxY4OGAbQpq
B5EwlxDF3Wor55CFE008CwugBy/jVMvOiXpS/oYRT/9gycWQVf8efBrA1EGB6E21UBqR3C+wuh+S
oxAbCU3NmjfchKEnqMQ0zkaIq/QwQ9juJ2Z8ASsiA69+zLjiYTX1dAH9Ryc/FPLLR/sSpSTHfu10
pl6z3duvCQ62xtyHVBfGkfR5Xc8EhWT0q/RbVYJ3JTZJN7PQuy+OWG1PjyQ9rnN2tuAZPCaNUI1v
8QJII150AQpzxtmXBqi3sl6ZH7nB8QbfRCtVeRwn+QsY24jatRd3dHUfbmaQmsD4S1eLusCRFZIE
Ed1Ve+8V3CuHk2CtazqJhs8yMnBSHZdcwF9A4U1bAoHndFPgY1er6qGUPH7FA2vds13291bGk3Hl
vEuc4ijDXvN0ufb9rTtkZ9ptzKxYOgqxOhYjaycQnOKXFylwWRtyvIL5jwzGQQnLR4lUtoXFn4Kt
v1Lf9cqu4Tl3AKqPJiVh5nGJOBo0LBG1h4uKVP2BfJGQrog0TGtFzf9YuBIMWA/MXMyOoI6Fncg3
BgfaaZ2IPNAIm2TXWaAly4upfGvhxiHo+KZ725cS9r8SmQXC4zJID33eMVcVg7xgjx99DXcpa8Py
c1GTil2LP7Illj5XgBL0FyAVBXYOGqg6k+13Y0NG/5vuGXVEGWZCJ8teDgLj55c2kzt3nHeAp5f5
iq6XsyoPXGVQ13FaN5EHTgRyhEjh+OcjuOMiE+ZgKQBQ6qrFowIxPneJO4370t9uBmrKihuqg5PG
j7HFV6sDy/n7dWJDUpXCugiG0dQV+Z0I6rq98gn+l+vvu0du0DkuhgCbVIGprMMG1bApCCqlP/34
B2dWIxDYvtnl2dyjO4KrQw6C9MJw7eRFT2cctNOBeO2/E9K/6C/ON5VbToAMGAO475+xo3CjgDkc
r98PkPcIJUa8bqfisgCe40ldLdLQ8ZTgHY+KQ0OrndM9lYhLOGDxSUk+K/mdGaTRRzuqSL3hf7wG
Gpvf95cuum5whxietPOzMeVa4lMIgMaHiJ3VPBwW1EJENvVOwMq+9KnGeAVXUSqpunMTX+3ZVmUy
XN1/tK8v+0GUN7eKTVvDf4CNr0cNKH4sf61uPLMxFZA/cDLhydjEs59Bh8ppYRXjt3BfvLJ8QeGM
+gCe0DUvdjlOD95lBSeV0+IetzC51ArzGyzyNVS485h27xTeK3mHZuS1z9l9Q57UKDsx+lsQcavE
vKQ9CpLmt8SpsYMQlRIWC8wQydkiIxmO75fqgnbzIUeamJHY214Pnh/dxAROCKcFviibU5iKIQGj
XWXG+DPk3WMKFtawFzZD0j4crYYwrUlqTtq8eipHnRzrQAqjnHv8v3pGDgLsBFKNN6XItFkN4BYy
HJsciExLoefRkoxbfu3gBdJ0hlr2GPOIqS59O+sTOsPJV7ziA0O0j+KCTYWAGjr7oUE7WvbLX7NI
3atbdXuskZ7Tjhqm7CcH+ptC9fHG9S4Q8cbTxsmud73ZoCnIlgpj9sWu7P+/AZhddsy3mx5ZwFiz
b01fpuK4CS1Au7OO+WvPc2jlbt7QF36+AdI8Css+g3FaRLtoG7hbP75opaLeKl4wJVXV06+yOBr2
lY+YMl+rtnINzcbpQJPeisXi6uQaqlIAKw/gkRPVuvyhEqGUvbW9uwzaOn5xvuB6GbASwKxdWKX1
qwpfyTpF4iRAqGsFk8Jd8sGD5xP3ZS1RDMalrm6VYJYxeCHGBtXPfsbyDKINNDgIzHJPA9CbgdTY
GFwrotBRH+hip4mExfs+sbyEuJxG5jwg8nZf6MEGPBBgVhdV2vcX5VYTIfcbxVhyaTeYKcak3bWl
r/mWNIlK99co50dPyTZJieH7eCWVvDrqR1eBTkV8HMubPQD+IDqgymdG9AdMNOeggDrRwGYypP+O
7lNZM815+0HwpT2g7ioe2sQiD41Bl2QvAiimI+RoO/n2sqn9mfbD5/GsVjxvZayye1m/kj3LtyE0
94PJh7uAkMzcj5E/YXy1UhXraaxz6X6Vdc3jTIiDfzmfjsML57ICxr7WQ4JtehhkgbsWrXz6WYtC
V4cp/UcAqQNWSXay1th6PEIiZeKIy0c1MlrdCXC8KBopk6F8RzSM1ZxGo5jrfa7GO+Quqh0ZYMsm
lZ8Noc7xpS4VxwGL9BornzQ+2o/an70K+615d/4xk8ajIWw4Fuq9vfAHb+qBTWlY6vdS6p5Q59FZ
dpUp9D6GmXSVm3eH7IzBBJ++B66uTIpJYJiyTVvl0fBMuWmvpZmzEUQxUB24CTtLy9vm2ImHs4Rr
dMzKQlI3uxQfPdGmyhY+v0LuiamCvn9eEbnYNhAwIV4FNjYgoboG9UydhnmWE9rY+qaA5T8zDDa6
7kzv/Axnnrtzty6/wKYy+1+nRlzmhH8/3VM7sBojRHbK3eL7LBb9pVCdwusUN1yD+3N5uemFcfIv
pRj8zsMwiwN1CE5ssOGpX13W4ZT6ez2s9awoh40VXVysBqBToDROq7t9TcagIZX89iWEr+l33jY8
sf8XxfEB/hHWx0Vy2jnqxcTIi6+xViOr6TjJzzZZhtvtWvFyKxnyQWdEzaovBQCL/N/c6B2oXMxW
jaVP8tefw3zGlSq4bncvl+OsVxvCKY0bGLljWPUt1bQS6IX3F6sDxYY43dHmN+aZcKNmkyB7/oxU
Zhrhvs9AvPs7AcDJJuCu+yb5qh0bOAWQx76DSApsmIRsAH2rGvTE7mbBkIWC63a2Rjm5cI/pcdQB
hMIr2/LWfmBGodjEiXDr6oybfyPBOwVj9aYl7dG0mOESEVkyimKh1zwBoxlZk1JadQgs6s3BvWzA
mP0u8jUjN2ETfGEP+5Wp2jbxrZCwR8vTd59rRUbd05tGtafG//pwWAGjE7MO/oXuiBvKlaAgtUGm
8i1MHCL248la/R90wHd8yZyJqcEQRESVQfe2epBaFoTRuTnH3BOnVYoF2PKmw6Dd9bAQ7AnwSVMn
rHufeBTYCkWkBgRoyjcxWtHmn9cwx+3V2mPHqPfj9VFiOpadKSSHoDYGgtctlJHBCfM0O+wmIt0R
qW/hH7z63qnWvDAuyrvHNIl7nWTC91gnmRzv3V4Tau1sFPJlZCuyryO8ujechhKJOpYhSIWe2J+H
Tjo1So8Lf1qKhU/UUNwk2tKYn+J4Y1tE9l36161cV5CnHManFWx4k3thaDCgtQHtnghqvpogts6B
iIn42csIQzBEQJFY2z29nO94nCxncUwHUIWeRerzOYPYMn5zGfvo4H0NmdyGvXygopHzthkSrNnN
JqTp5ge3QGxoH+RznTM/+paPJAIFHsBIKd11VG68eu3BWe1f802cwcMRZJIUvObBZXW1EWZRHRjp
SuOM7otdTxBIXhsxNAaHtHN+7FbcS8Lnwn8S9kfqxdaFP6S1K/7jeAmrjn3luV7hVPgNJA9Jnz4r
sL0/DvOJrq4SFRdtTgXTzg8yeE5+byd9E0D4ciKp9vaTs1UQrOMC6uHE/7pTKdClzuwSIc6we3fB
DhkG5NNE2posaebOLhMg+T3l6/svWaW0WIffWpKu66RDwceLAFTCVU6zarUKM3Wnnpz2PK7JhWey
Oshahsnsv0ahlITH704jKvI+GHBI2MvBkZFes/o/uXOFS0GF7Z21iYLXiLEhEslguQ3H6mG1LcM9
r377EE6COtNdNZTf281TawDKE/TyQ40SVI9BNWCp3EknD3Z26OFSnd2pVY4olWNuJrThsT4MwzCv
z2QACBf1BQYi4PZoU7yO4pvxcoS9kvsLMC0d4x2UPY52zb+kCIXHZ6EB3mekjK71WEwLkGgXvZRX
QOJWWglk++96zKTxEbs6FA1TfvDoxf0gF/m4oy4Boo4P3rFBFZ2aLamgeGnXzdI/MZFBA9++tdED
r+qiYwPeYoKNpDoRlF3kPS+8vfnjD/4difAGHqHcGscT3uowSAoloHWcTBxDNr35XeyHN2lO9JMq
ix2BBUeJJIjk0ofrdE9rxrPFRn1Y2o/e7i/ART/LKGRxjjTwlBq/2pZ3/T3Y1c8mVUKaP4t80Gjq
FAWXMBa1tJwbWK0gGsc+zkpBAQXRZfcIPSSU/D1809yS84dC/bqvZqokYZvy90dwJrABYOdHKN6r
p9PjSwiVuc3vH8l6PpTZlsyT/bzasfK+y9PfOAOxwHLzvfweS+gCqvKkNa6nWRLH8j/xu3e7Ngcy
SLHKqFLmK+C8FB//ZNojOOfAeAD2iWlggXHdDJ759fSezqfnx9n2JxbH3z+GIThhHKZzw4tsG6vi
spmDo8Zfunxz1EYdMwhrNEwZKPIm0Yr6cm9C98axvxOuZDx5JKLa6fQ0FDpQujgJdw76Q9qmIpPF
Ox9FVA3Ttkd3DylFDkfh1ev/Eln1ULEniX6fo/BIqt2pqQaVoeT4id7oeRj+PV088hk6E49BpX60
XmYozit10En7Pxulh2JVsgZndwyqHIaXqHz5qp7a3QDODaOTg3O8mi9UjKx+2mxpHVOEE8BU6h3r
sZBnCU1AOEoq9vp09kicG/hmlAPP+6Zw38EPyYfz8A79aZGe7a3UyJd7gLiikU2g1bHhGf4P7zQ6
WzjAN31o+EvQYAwg/LYT3m+aN80/iA1S98CnaYXVMjTvoYEyFHTQATv3iNW0cbP1UoNtZZD22nId
cNZVKRw0fTu8to2T0NcBOG93nXBpDIkKGoG9znt/UNuDf5ZLyRt94Rf54E8FJYLjO9chfAtR9m05
gxHVrBllljTVmx9Yk2RZkTB1fGShKUZFayJQc5e6SB9XQ10DeXm53o54UNHuZCcEppGqvWY9eEoU
Jc65QpdC78pk3EDTXHd4S/c6oF/fpKO67mQq14MjtTnvn/1NN/QYaSRoJdAF9X4WeQzAZsXB5eik
3gKrQoGuhFFp+nw0xy2YRJD+2djW6jWu7rvlORVuqv99Jd8tAv1QBdBt7O239dpRyGTvXTbhmC5p
yMORK/Rpi+nhmxZtCwqmpeWrTnhB/HBuK2roTTyXoN2g4+UPaXs3cw7asgR3AKeK6WCZuXi9Vs3h
A5T5A1bWoYE5I+UDo84WwbIsIu0xQjJmig+fHZridTJqpKJIoLCOPXv4ooNvIZI0OyiiaAu920O4
rBTsuGd6GigTtavSjoi71qDLjKzkc934HDeu0m4/ZTdn78iIIJ5lHMKjDWmAxVtBxHXpPys++A61
86r8ZbkgQLaSjA7jMt3EYpsjMvB+ivVIFUNNWu7iwiO/i+bb9KJiaZESu5YMzeY5vlxIC1hZxHmk
dwKWVk3rddTAHHRzSl4ddvRBZee3vMo5WsZiiMCXWGhvOEavloJIik4Q682Db2ZBdiRvuyZSG+DK
j53dVyUPqfl5zv7Hh9O16yGLoR3hGnF2AP8dnBgb5O+GbCzcW5ZeqCddLbaso2fRMT4SuB1VOjo3
CtWMRv/18MejOAfIJVckmPijt0+bwuzwagWknhc7YBOCeuMPskLDI3ncSK+J4tYUTmyjs+jVrMUp
uHZl2dBsuUaY1BSAcVFq/myHrHWpq7LbItrVXd9L90sDWIobbXooDkSG2H0085KOZkLl8NPJJtwX
8uT+e8avQqor9IeU3xcLoTO0gMghAleFHGcbD8DnTk1ieISt+Wthv0pjJw4z68j4+exNYn2oSwvE
LyLWXBGdoNRmdew68WaJfsK5YXcF3XnX4yIBZqTAbIDAdnf7lr5lhqu3Kqix+rbaSeEJvYsAt4dz
MPry6mQl6fQsHx2FRVoAMBSS9z/DTdNMDchY7KcHDo+LThl7i/3uDnVPXeLv2KBqSogF6e8qRGUF
5Gl5g+Jz+s+PUEAoOKuCn6OSoOpujrGjTL3+xDhoNNq78qWKNYH3sg0nDjMSTf0HjRLs2W/uq4Qy
5KDQY1F0cdtOhOnIBXIHEcdeDE0k+ucTY9WIRaUTXmJwxRGratHxi8L1IsdKNttIROVp+Jy2YyIa
WzQEsKLATercZq3mGmL77wyWIAjvQF3ql786l+/YRGkDzYNc7u/J0le2g8trALzhV+qo8uHu7UKo
6GcPxpI/xKfzKU9sjBiIUpvVJ5p2Bn1qNuZJVCITQcJCrX3cW95e19+dwfox6aUzwYcZc4fKyaGx
NTos6XaWIZ6qYY3ZcIlkJjsdPiFiXTvMEcNzYD7i2ePxW9SiNMN6fbbMe9P+QbYqObGRpsZ/oBjX
hZNi4aJtvKtb0TKRjOzerZhU2K8/amBmgb+NhlMCUixUpOpypvcKH2CD0+GM0Zfc1owYVA8Nxa1/
mW0Lt2uX8VkaxZj+shSQQUMmAYiiVYU/2tz38ypmRDPeQ77NKx3SUC0IMC93yiQMrPxOQaHjqXAJ
v3gO5yyOQjiUdslQnmLqamrQtxSv7W6jORh3rL7rYeG2Y++Q54rRUnhSjqjwCXOCDb6c9N2vhP9x
V2IENbnFu5e8Qjbe5Zbhys1fWwUcEhs3dMVbp3Tn5hYGswmw1GS14OHcnp33RuMzpVKKaFmMfO3G
/YXluo/GgWYu2wnJFvVe/EBSSSdJC4jcdv7ozeS0Dom9/YMzvrcvwgc0VZcFRLo4+FcnajjNSRXS
Zb+2XdAUs6TYn3zTWBEtHJUP6awKPVgjWOtIO+5UjDRibuBHRgq6WgveKqUBPFtQZsGONb48nP+6
LWdb5lGl1GfNLyK3UwRrBKM7P4IQ2rZXgClluABSmCstcdBOAWnBYnJTkG1Sx1h4+9toX65WIzsL
FY0BSl+ToGG5jzW7Lzm/5/FBuKtmg+KfCSXN0KGW9FSwip9OMMxKBRqH6ykcRMRbr60bZw2tcrMR
mjtMGrcXDLkkMxB7TeeJQOk1sIfWxhQJyCklfrykAC0lyhzNGQ+IDmaWYjbTf1cjmXXCw2I6F/6m
CMldXx+0e1r/GRtj5K3f2lMwyruebqKYgy5FiJRuiNU7Lk0uEazJDHiQDWLrX6ooMpz8HPlGdDKK
mo1R/kELqlW+4V8/Ca3zN6fJEK7xScHxYEyCh9KLCujCoXLGM2u8jto6x5DZYycI2N1rwBrWG+Lr
FQSWwjrmKLLotpCVwiik5uuORFw0NiynIh2tDvp3jPCCeWiGE3hxzY37RCxxIIbwflT89+NAXDZX
mEI5X62hNUoXMCUyWYcwL3qbWX0H/q53EeXjxEP7riAhlz6Tr9mQxcRBJQHC/QbHbXtBFKtoaW4X
elPAngN0+J+HmssRRw87psiHiEQtSBQJzCuNlQ2ysAyZb0e15PSq8rED8c4xSS7fzW0fvbL36bDl
M5vloigy27lb9B0aeixmmicW2JsSjFA1jEEEy5y2ftwW1wlddPBsP6MNQ3QsFCXvdKiavF8d4kqL
GOqQqLG82ikwwn0H24AVL3upetVUFFnTgyGooYtLhpQ++dUdj+qAxgXtso2oJgt5IDRtm8Qw5N9M
KEpaczqvMEEJJpdqs2RsBJBAaUW2N7nYenIJxj5fttjTyJBOZsNL7x2xEQ00ToKJHcItXVwP0ye3
DI67LYUOYw025cwk+UKENGPl3b+oFAb/JDa2BK4wa+1wN3XaT4h31PrrnqSmMay2pGjbvY3KhqyM
d4GgCBSLPo4thX1Zbnl/OXjG1XOGhrjdU1jQTtRZ0CUVwZW71+NA5zpoqNZvnPbfEis3AKyROFsQ
Cm22KoNoWt3oBv7tZu1dZmMSke1MB1dcEjQYZOVCGG3ewyqodF1ry6YwnBojqXLmYDLIs781u1Iv
5mazIIQRAr7sbfzTsc1qlCVl7Obogzv9UVU2eqm8pvF+0TtjQWY0RaF4bpc7opAZVVkdbgi8+3zU
OCYIl+vKRzV2O++4GGQXd4q8vTKeVm9+Ko69Ir9pK5FbODPhpqfGPDVLHyZ+UeXzb/UQPPEG1uHB
otpehqllgxb+jLFBGOq4vC3iYDmJslqOFuQXNMtziEo7hIFD38c/xEyJTEmBLrNHCGy54SYwAe3F
vTVCXU3iN2FXuLALZOTJ/go1dgKmItEPZr7gSxG7i9cpSH9t64n0mKQO0WQuflR9mh9gZa2UKaKA
XxZvKLB98yTcPR9zBOZrb3BC695uYDssnj7sl6yPp2rF+cOe92E03hWIspMrtW18UgEv2XY4RRli
U671DqaxoAexQmJEZ/FIfqJVr0uwCGG2c7YRio69gksgG3r4mCXSizyCo4DsoXRnUEoYjCxxK8jS
kO1aClh4QhrBzbq5gP8YxG9LQsh7rfwurQjkv8EyPXPUiPLmMaFkCU6bNCeH1QSPfGjjz8wnaaPN
Xk6V1iwvjOYyvsMmqPxLSO2AYkcTcstR8E0HcPkYMh8RypidmzyVK3wRn4T57i7Wu2gqkr+1Lz/0
NQvzt9d6bYFYT2tgfHqHs0W2J0gmF6GA7HlhiJV8wKIKDBBUTjH0d1GrwhqelPpl7/afKYMSuI+j
OYaiz6s7ixaCxk4Q9AqWdozzoXYqzU4CGcnJc5H+P3I4fVhDV9iicFyEUmQXzmE7QTQV1jq70fhW
CATqOZB+QWBkjEl8rZQzRpXBqL7UfInudoyeitM3E0oEgYc/8edePGrC6+h3RXcm3OkEON8q1TDu
e9LKXAbfBCvdAVdv/MF9AIPAW5DTpBHNToPSrh+cdaGmUZLbjFy1ztJslzmPQ7LR8hPui+1XxdtZ
TjCbehkcb6N+E3AnPfIMGK7kbSQWB4aZGXVfSUepv2IFfY8UlZ3MI3aoDC7ziG1SRejiMyUREVLW
h7Uot44PF6/xjDInaAsP43nUJfguoFSDZPyHRNlYln3jHwfQhtoi55Ir65vmK1EC4Qa7TJ16og9r
BpV7iD4Pa1pbMNvIxFJNLa5RV0N6fdB8iUhIvOcSC0fWBpNpktYRQV8VFA2QOdiLYQOKOewzwqL8
05T/KW4Aq+gtIthWbiS/Dm1QAp9F0Pn/+pK7k9dEUSosZp/03VxZWFnxLpHREE4/TL/TeZzSpZIl
1czbt/vnrVUmzJmncHT6M/Kr/D+P43wYTmIItL9kghYFtgfUpT6wFfATueL/PGznI87r/LojGDKA
VkuVea5kVD+3G9xSRg2nNjYvk+slOlX4ruEFo7GFpfPWI8zpqylDAwWJSEzFVfNarNKzgo/WnISq
eQ+7asU+AfIw0+0vhxzheCOcetNT3TL/r/rFY3cH2HLYPQ5a+EooHV1kD46+HQcvAZf8AqMpJUKq
dUgAQi5Ho6dYn/FFHPvIqhbqx/nCkYFjXs20U5KRHLSu5OvWZ01G/fM01TMCiTv2Venwo1acSV2O
FchkqD8CHN5JWtx7Nvf1JiZMbQrRKWpWRhY8e7NenzLp6yjt9yoWi2AESDKt43ubTIuIHSaNltAK
pM23HhbXjqx8ARE03tGpgDh1Tn3FwKVd7SvywIMAGg/+jhVvaUK2JOGxcXj+jVHpn6GXGCs+Vrn2
SNcRfxAVI+geG4ZvFPDqV+lMXLfNSfUrVb4dr5ZjXxRh0AXOcyVm8r/3g2q6EMiqWbF2P9IDuPqB
wptJodAVWV54i9JImT5/o7XhMZ9PLZPdO2iUEsTRh9ykruhJiUrNGAuKi6T2v4aVDg5e/dYii48+
vCToSxx1kPSgm7aI5INvM74g8blQC2glUsy0Pabe1Y4lZBF9SvHT57uSMTwzbvwjGoWuyEZxoQlh
jG8n0GAtxGAHf6C1+35oVZAbl7oOwnouK4V4Nfw8ZeyWQ/3mPOmRQXMWPT8r6yapsb4dawZ41CKe
wxKscpxZPIIXFeq7j0BI3XK7dYkLw9W2Zou/Ipit4eGO5xO8kt7GoV2AsNaVDR34B04P4puNBSNG
bT+aLghwJbmoJXi6v4Os6+0qHHM+Ca4JDVLZQe61BWWg0tTrzi/poaA4LzwH2zBpe/lIY0Mz3l9K
FKCwimCybboA1jJtDyW9P7mtJZEP/HD7uRGdNn/4F6P4TyYTTdTsuIlOrnYU3XCEHTzly0B/Xe2w
XrLVSXNXtOiaYKyV7mFiYEmsvDgFPKuVWtm9y1GE64cNhDRe9m9oRLh4AgUG6smaB4L5p4qX438k
Udvwe7EVCp8Q8d+Fr4/BBVJwakDiICHmUnRNZKokt9d+/LEIQmi0Ta4uyoB3YJwcvICBUJCO6eZH
noyu4sc1dRTa6c1z56F1rknljO65oihOsFg4mgmVopR5apmlZdOa1WKD47wuveINtCALv/W3xl7N
apI6wnGLCDPKrFySmEmD0CXuOGBI7hK9evTp3u4fiugnXxlYWTVquMybn6ARyW9Y4WcaDb+mhvA0
T9xB163YYQSFH92UfzdUZeu8knKVwIDCyxm961zr9hlWLmHwhcUnUw5F8lnGI8fjy0RGojR9SeMk
FbcuHejfPO7gI2Nn2Yk9pnO6criZtab/wUZxjYtcH4k9vn9dcnrT3LYi7TBx7fyXJeIQN6GCWNkA
/VifEPuwDLGUPU9pd0D3DLdeiRxdHEbXo2mX//9cX7Jz8aHwPdC/LC0jI/t8DnzFOQrXb3zjIhjS
cP5xqzkC8hiUBMwj2r4xFP5xfqud38nEmcVBgkIJDWCgE1aM2tYQpy8G3ecaRFMyv5i/ItS2L7wL
Gp5jt98y/1LemybQhwTIaZgDZzenV5cqewmZktPXzG604/l4NpR0wZfvsAxiHeaPUnays6f9YhB6
dJM+WlsegaEVaNGfFEXEvYqOMyIpTD0DBQt1UtF+PSVC6EJA4VCxFiGoeWXwfnKjEJ9UTymYLNkN
gGpqxleKIrmcxDayJzsI+2DvyZopTMM7e5KFRkVP4r72F3FXE3plOTvqpAI/6Xmvn1danT084rMH
wEKSYjgohuhfySDlt3bxgGvq8VKHsmZXj8pmWANRqF2114QTLHl4sYGbZEq1GRn5z24ul3HcHrtc
MILs7NIyjwzczpyphrHi38IbU8p2yRM13BQoishIKsFZ1G0pLA58+/qYMMjC3k7hhYxWTdDRaaPI
amLTwrCEZX1XhhJ++WZoc30pm62UAYpECU3lQNJr27D4GM6jbWlja9VaEdjvnDrthqUHdZF727p8
hGmbMHRWJ06yJbpJ3JtoNFxKY3XwTUZ1/oY7y0sq7SYFXnOoA7xs55LFhDyHoDFN8GbUnmTJqPft
pLQ65oqRe9NDcwI4PRqLfvFw26Q2QnbnR8tMiHegYSwtt2VM1BQi5Ij5Xj97Zecl+gbbgTg7gLVj
1LrciHruK6sGxEN4mZKeeJ+2CBa55VZ2+6ax7sSGAXL2UGFmKSMu6KWDTclhk9stEd3kSw6w573Y
GF2pukYA7JQsDQ4W10BxgcZPkyK6BrkmJyl/ufIvJHuGBr5koMEx84J/2NnSdIY4I8BXRbVJ01ZR
M5Trp+aNFhPGFfmeIhcMjtNyPlrY3QwvRu5q5mOiFWAfT6Gdlf2naGrG5H612X4cc6mNp6YaO+ee
jPn16K8G2h3hn79xZXtNCERNqH+QCNkrzHlQ9O0EqOx2GlKXKs6hpYy2nmdbzk6o92qKoCBaeIqE
4NeNugvy8mudIkyw5QEZxeibQaYKcKglfX1tLQ95F8TiWfZJJnjg5MSEeik6ootHmGKgT4iNo6iq
FDyugP24Nzy+NA3Q19TTjs1XUWaY7YY4+teuMwmHfyYp80KFsjF0t5Oiseww81oB7gr+2V7LLIck
AzcTo+DegXjYj/96EBaU3pawxrUih5oZR4ZezoAeS+Apwx7tQ69l0GIF4P3s0L+98OHF9BoTT6nm
qWyzEwaZnyfllRRxtotfXaOkAkDhmpuy5JcoQZJbfzM6NiW5jgu4BijQvrQd9reol8p1OHv0Cxdv
72sPWgwASCax2LguJS1V3a/QtL82Cn3fNiBXi/ro5cZd+cr3zJ8j+vOXPKkXkwHYJq95uRn3MQT8
CLQfAZL7coBO3480GqspC1y+NRB2q8XqKPmYrvY06khJEgcSsU+jPGyXcj84kegX6A6lzc9c9fcZ
38fsXHpDQNHPf82tRCsNS403AvIzxSNL4QIHeNBlVsxNvrGSagoM1cmZDnBgHy3pKyjyXw11J/pU
dq1/3FLkhYEot8oXdwDeNVffwWmyLoGRz+8oBA0SC9f+jFKkh3w082RTWOOMo3PPJeNMX77WIisJ
Q17qwA/pyLqbi1XB83wyxHoONVyY6CBX6RhJUYYMSFoPak8jfK3Pxd2l/e0ewHNEeJMdx9pRMqHt
Go3JuACCEUS6amjl0YBOea1DUMBwMaUIqhRlW97lMwcx5z+WZLcgvZnCXFw4UHsj12rSLtFvGxVl
NZzVaIylSq0KFPQXKsBxH4rq6jIGlp+xgYYw3SJu6bopaI0F3GbeOP9M37S79xG5DB9w4pOFXETL
TgulA3nfid1wlU+35DalFFaIbS09Z9gbOdb1tZ4HYr8mbIqnrJB/aXNov9xsi6GQTtXWzdQ4anjy
KUU0tTSsCLkq8tgq3Ye1+LwywJp1PGb/YoXn9eS/3liMxugonOndWRQqogSq6TjyvVzTphu4WQ9h
/KfVG0V9WvLryxmdZyKeZtp52LWKiQOrPk42C41fPdCEsMbi1W0fOf06KPqaG2DsHWF8GCopVhbt
lMNOO7DLv+1xFSCww+E1l6gpF/ZPP7odGtov/2S1Z4qwNtE7zDLRPQw/LipCT2YnwWxeOCTQtRfH
YFsMGVVtSzxYyV4GzzygKJWIjBobdrI2SV+ZE+DmsHhqNEFBFZQkFfE1s7FQ6hHk9abjGwQ2ZBl2
7hbmEZeKdpDd5U+Z6Ee2hHZKX+tI/DVXi5YHUmNAocRoKLN5m5nnHnZJ4upyPUg8fcy91zjlsxzI
reMnaKxoY52zbptRyN765qz/IqBJleWRZBXghhka0/EvlyEMTlRkJnNY2s8YN+ZWEKC5qMloSoUA
B2GUdvSKBCXhUt8F6uUYWx+Ayfd2rAYra2pOm7ZsJb593oRUJyvCcI47QRbs8uMpO4kDoxKKUs/R
+dMxaZZKJY/FgRVEuWFeOpOFI8cRptz4eS0BvBDqOG5etVFZa/LBMY+WZNZGgcfDyTBFc+Dod55O
7yjTz8/cIm3cumvfys9ZKa7fHTStcK28KGl5iTcYDLIZlG0K7thtMvI+35Ryz74fXzv8PAQ+Ex61
K3JYvkipmTSlP7S8h9IiZeIvRmmJyyzYWIf+Nui6bt/8T0GfaDipbFOcRlRvx6efHg54kNvkRz7M
njHvc0X5RVJdCWk1IZN2UbIXPFvbQrrofvFvKJNsEJR6YFBlrf5ttexdicy0RSYoI8X1S/X1AhDh
gtokylk6Wno14Z1mBRLbb5kvb5hoS1Ck1HJYkFZFO8J9q7ulw13SPOjply29cBF+eSmGj9Mmhmqc
NbpBZITqyk/0acZIEJ5htdTh4GKQnbdaMKBCXu3CqNmivVFFFJaTK5q32IoAzr4Zvmen+zY9rvu1
MBdeY0ZRWjTcmIZ1v0jqHrwzpLndYXVMV3g+CY/JkG/orVqKERJVGu3mxhqgz4xBBkfhQkbhy12k
ouro61f8OoYW/wcieaJ1hJGLtaRkTw2JxaQ3XeD2yltnvMXPi7NYraskQ7sHmx8gnB5EPEziTNiO
2j/UO+XZ82nCeTlP7HCEm86gxnrhVSG5e2EFdY0DRbrs2ACEgr/JOalv28LJcMtI1RDt1tNyhTU1
FeNSHmZga2dGlvs0yIoACCWPr7WPn99WhrwH6Gw40TD8vWnMBOCYDENKbU0kZE+TvYtCfnqEef9+
8ZyoUPaEda593ivqdB3ApzPSGJkVgjE5Ky7sptVW8RkGAYzJtvPgfdtQOOtUGidsDaTEOC1G+B62
WS1b8Qv678AXeZ+S/6dmpJ5H1tFWTGd8vThkoMwq+J+Po4ImKL/+5LYPVOKWkssOUtkBud/Tsi2L
ZNEmxq/hXv3URlsQWNMSN88FrWjwIC6qymXQIta+uyFCug6PSmB3/v3TxamhH0sDr1njtUhB4asA
CMrCq02FjAfv6UWFvUSrvhbTljJDRiZzAdNEctak2We3rxx/mwtbxFemh1mdCrkly+mj1q6BNlP7
OLGfkgClG3koH3mdT5vrH2mKhvgdJ0KyzJu4pL6sN8NtSXaSuuv5Y61FoglGpTMpT0YoXOIBhcRk
Z2BXsklMlDFEb7EHYHbhRt/ihgiWpHQf1DzgErYbV3ASV3nk1+jpqDfn+QVRL9F+mZ6wWyIBTLJB
K84uJmAc8L0L0xxVk7zpq70hy8tX9NK+rWM9Gn+6h9nu4QS3mNlk754czTusOMODs/ikNCfibCEd
XS/as99sfLQBu1Qjvs9OqMcln1fi0Tkwh55l5uHM/+siZDjVs0hUJYwWyg31uX8PLJ9v+eLa2bQT
nmRZS58f4WiXqRvTeZ+X177LqNyyYtOYFi0vGkBwFGPt1dYLRzqHwqSxPavtnMe0BcfyWMufQ/AC
WdKDy2rxwhCF5qlRvay0EoqYR6EoVvyqvaSNRd9ePb03Bz3KvnFvUgmlkDuP8ILaapLikHS3u0zp
zt4poustmHzL4jzfx/57kdeVoF0gN/bjTS8OZcYvRgemjcTY+Anc9c6R0axK31e00/euTe6dw8ym
c+IeojAbYn26N5g/D3OzxWDNLiXVmZD0CnRPhuv0Sj/uB2CQwvGVR3qzfmu0vTyMe4HOwLRNt1Qv
L2za+A06CdP1zhSISnmHIOI2so0R+R3fm0VPqfTR67Z/iqiRZkVEAPPkD0hJFDl3+wduBO1jTEL/
QdX6GqYfV/STECnMQWLdslwmBWTBUJ1Ixfd09tLY/ARHhEMc8ETrOVNvDrn4U8rx8Y/+q4XQNCMZ
CC+lwSjxW3hTZCMSvX4muKk435qy3aGeKOZe2u9SQmwG5+lhBnhLkDLvTzUQXYNc+VMyrj8OOccQ
7PI820xiEeUJxnQjPFoqGliKBqmJlADVUjszqQ/zq/4RT4lhaQQYIHWsTe+g79EIHP0ad9CCzMAB
ljfKDH5H0bl6ucuhWXGVuxyCQpmD2/Mr9axOcSPiObgrhTKKyhN6E8zt1p+4hrONvUS9v2GjFLOC
E6zFFlZiATx314+7v2r4pa5UsMAimKHwr8XpZTu9pPYfJ5qvtkWrbZ94l0JEFNsokg5rpbHjM6Ca
F24wPNtNU7hk3FOio+QrPsn6rnf5na22PrAw/P+W74JAx/Xy760RYaAPVVorTR2oTd3gIefnWqhb
+vFdAwmoLu/Bvk+ZF2bbDokDMM50Pgwt1OuimyalMvBVEoWv5HdB+CQUZ0oRx2x2sxHF1aejtaqr
LEB0AIuS8wSLRrC/2/ey4jVYldPp9T/ONfD3j8/TdJ4M8RS1wWUunZrTWKs4G3uiHhsHocZZBd1Y
olgdnucB0jUmOF80+w4KLGnqBl1ETj/yfdOt/L7scob/QAalBtUjMMBEZ1hKbmnLT86bUFjN0FW3
PKxLBWTt89RSmGYeOasXVyZeQ45mluc3+EWYWY6MSCLURUIUb+TPHKea0jh7Vvt24uRQ3wv1Wrtv
nVFiDUDcZKs76PxiJvahdfz4Z8Q2aF0GDgmcyNkSiOGX0j4wSSVIUaaubUiniRvmsBdkAh+zS51D
lv/JTKbXWXYNVtiCEzGyn7+pWwceLi/Mpv3d8zHZvyLfIxkQOt2hWQ4g3EH90D0L6/dZTYQFtOn7
0lHZhb+L3pJ7M1LOH1Dkb6XHxWulJ7SKczNJvyPZg5H3gpyxIe3vg9e+cyaYx8g2RnKgKwjUfn84
bX2A2+u3EuYHuItz0/tf3QNp3B6edUXMDHvuoJufy527Hs5HmZA6OmxsOXkTzosABGgZE3FiKXRd
MjwuPAhwnFuZAVX5fXgOXiQkUYcJRNV/zxAlthC1c5i4Bg+QWGfCVakcDrJjJ94lV5bI/wqCWkA7
a72IDrrmzl1Zw5oV9Y8qa06NnYK3v0istefMYkazaFFVm1VTydq2flf5meftHXDRJy+hWl7YSaGS
sar7vG78Q/Xg7VzNRZUafq2KQD9aVpKjLq+OsvwPhi22Fmygtggzf0lt4NihXUrmN5q7iI5ORuWS
ZMG4apE/SpIX4yYXlhcu8lDI6MS3n14FvKMd42/tRRNKMUB2yQJ8gA88UmmAaQC1vI9Ljwh6A4im
tIfdeECDiPJpUoGEmf27LcKDIFrKrKvgAzGmRsNsShafcF+T0bMcHuEyQa9OZOPIlzdXQPnvI6yC
B6nEb7ni7NWyldt/NXwvQt3UQ5KS8v7TlZ/FuZhFnB7gn1BUMdlL80ZnYJXUItU7H5lr6xX4LgrP
U7reMUj42CvJw3OXkmcwLh07ojsFPQzw3JItk6yH+EZ7yHy1b8uK+lgfkbok/TrK8R51zmL+e8zY
uLjPGpobJQFFUNobaT4E2jSj6DVAFgV3bjmdXY5VtdnzT6H1JuigfTHR1m/nVyD5qii7JH12G4kf
WeJWY/o6azdouovtS2rnxx+wcVxqud4IAyrzdw2kcKsrFW2JDDzKuzPOyUuCttyB9AUM7e95xyQG
HVoOOhPVY2EywVz/aTN1yF7RbkcqSrqkJO2BCZz5OrmbbCMxcu8ExxSM4kt/43sp7U7Vtm/rwLQz
NXhaBoQRtz+kGmVeRZbiBf9Eauz6SNrQ68OFJ8ZoUeYYY6Ao0CXSOlO0qFmlXmpJYRQWbsBjT+9O
EO7JxUAnET8loZA4gHLpmX0O/akWj+6GLFw07f1eSkMSfgt3jni+5lYkP7+UJ/VTUxix7CNpFBz3
TTGrw43/ehFuD/KhA3xlK3/c/JQqIJn6zx93LWkQFgCsssj+1sO75GPbLYyDZE9Wl5LLnuyQm5Uz
VCs1rRmAXVIL4gdRsoztWuBn1VJlFI5mJN6deDFE56zjLkEJP94gstTSeVqUinHkwzIZuCWmgiqs
ZHCxnZHsaVVqYZfSUbficjQw+6eQQfqG3VL8Km71JsTmBFlOrjdsdKCzkmdA1EJq3gSQPcch91PW
dvusWo0cHKIE2GbleOl3MLX07kTfGvs/yc5h7EeIAKLAhUMWwAXlFZ20sFBRsCEesLsJtGc1yDyC
N91a3a+0UerVqk4mdY8q5zsz4FGLykSFjMUJA8hsxOlkLZsSUAdgnY+z9bcEbKUpygA2EnqC5Wh8
NtfN2SpIjbnv8lx4fearDw7AE5DehDlLn8PkWa/5t/zQHzmtWSEx2W8hGyBYoscnCTR13fV6eCy2
t6Hx6f664/ecWyw62F/oVR1uSo1pwNArydRD8BA/Hfsd2zarKteRNCZQfTYcvoD73kgZHt2kvNDx
6EJGZf8LiiLhFLr/yWxLtdpUjNYZiLNbrxV66LVK2K8dH8IxI9WUStEeCDVxGL6v2qvkduqsMqjr
u+6wQIttCjYZVDP/Fg+aqx8llaXcloz4n5zA4ZdSRvX1kBALy9dtjT4Xe13jTy57wrjhKem1l5k3
4Cjwnmhr2yZ94MGabszQ04qxbCsEPjv+YkyPlW9vNvp+yrIZrnqjE/y+Q3ho+FBvjiOcmSJNH6Sw
Ks/bMa24VWnRslN703hm0DJk72lGWo6B0A+GeW49KorFczNG1tV5iH3/daBRFW5BSa5SRTOl/glo
HPxkmuNsaBpmZXcZMOyxSPKcEjzwdDZWA9gE2j8Gcpo/5a1Kx+0/3fjBwMwUyh08PSTwE5tmbXSI
tsKltHzrM+LdActAQjVLGx6B0u8lumYoL8Z0RH9V12b3RJ2sq0nuU8GvRUHDs7BbYT/UBVMljjyw
Y1Cdm+/Y/p6SQtHQh6t7WwHWg8n8gnbdyGnDgUwE2uwVVfoR/jdrqaVKHiwFI8gsJsbbiedWNBrI
4e750fvlaRiaGsIx/I0rQwZ1oBBT27XAs90+FMs9iK9bsFOOLKLI5LMaeOXulWL+3BmOwPw1RZf7
PTxbyPe8uSu6N8EjEeRs7Mo9ml/y9IYOE6fJup8tXeMF3Gb70MnFbMk0UXD6lf2XucLU7sUK30ZA
xPsXtMEtHZtbZ+lJ5bxf4hfRFL1m3ZROzEwDYB7/UFkTP8fJvQaqaNgP5RVZuHYXxuv/XpdETglV
zOT2JHW4m5qdUajrOl9hFiiinaNJsQM/WceJ2NOvEK1na5fAP2BUfbVuF1FKaIJUoLC+2Uw9+XSQ
DdePGtkw9H7yYNpdaKe7sC4L61LkgyxkDYPI5MLNmE9mJ9DPqpFvBIOO9ZNuxK13EnjwZ2pdtMX6
AW3mp0KtIL5a8op6F/jjWbALmQyp26QtIL/NtyO7JKxSycuN5WjFHBgW+ipDIi+zl+mdMRf8V9zR
0ZAya1oTR8rypVidqYA2oALeZvchLf+3V6fpSO42XSmxLuk/O4Wdb5SXTAeBgP/6O44LOQwS1YcQ
DKVOtGyGzpOWhpJfgmPfj67Ig8Bq5RwGm14XOoOxrNHbRxhk8S0drk+JwAZmkCIYkJMobwSR16D4
sCoJUQrHI1+RzWVFTbhJUQeemlnAL6QcXCipXEeNSMHaFkos6frWSQVbdKZKE65vienIUykSGz1T
49vJDxvOMPS04ATmLpwFWKGt+3W1HESN4h8OJos7XM8CbP/0TbaDE0AeexyeP3qH2WHyPykt3naF
09MPWv1la1PxycgB22IogtnfmOKygUjQx+6hkpwJ9q3mqMFzpajqENqQgA06Aw1vLSLZChUZYFYZ
lRz7/c1vFpN+otC/SxN8OGDrwUZqksKSfBEvejPw/vbxaqovqpBsKCy75Y71BKUua9FsEeS40TyZ
kP1hbIn+a8dLSrsS2ThHr/8dbO079c6B6ltZa2ZgkpT9VHtroPH/pKxLIJ6CMuwSWW5+htsBCZTI
XK8E/FtmP0RMFAWFDWTLTn5d/gchuuo9Kw1n1H6GB7Bd+PDBcHbzyVJ7ZYUDmffRgHSIYvWvcKvv
ykeIXpK8l7DIBjP2kbMRrJfNidgn/L9xyvBDjcSQN12inrpuHwaueQbLwDU3fJO6f2VhX06wD4mx
+x8Ix4OHjJEebZFESlgeuexcXcRsN+yA5eEjULGnKBWqYCrSEsWUT4sFirKMfPYFebM6ToL3hC3a
MexLoVDAh5rYiQNpImuawwlANfGDJbBsGRsDuEfoG5tsoUYN7J/RBSOG34qd9qcj3zXV6CPWE0Ig
Xa6StmcwG6gMEE0/oJQWgXpaXlCOUfNPSahEQGLOhf3jNUrekgDND+3m6FepQPAcHD21fIvhRqNC
74zwpTez1l/nDDf6MPRkhYPiiuKoNJgbMdCKuT99S9zEOd71A50jPyKkDud3QeRNwXUEdQeaJma0
5hIVcgx29iUc2IBk6KiIvImNdIwt+3Ih/TKte/TqOa5UAolzKRWeHORsIwoO5GWEkKroLzMb1+30
ridO0qy+AKapLhbQotZfV4isbKzY+PyfD3aVua8VezbZWln1xfFtoZ6hH9vMREYoTEGx4o7BYH9b
zYftXZj7q5B18mRm9wyWDyuBEGZbRqrmKdji7j5hOCTjWjKD2mNj1ocUIj5XveiYhrB8WJ97DcU+
IBG34rDW8d/Sh6bvGigRjtMKkgILpFVT4hguPuuz9rGu0HFu4WdBmxJ7X/jZcE4D2Wt3ik8oHXfs
D9unKhz0p8PsoigESOz3xE+p21gourIG3NEdsJlE9MnOd1B50HsuWSNDgt2i55VyqarH/ELY5EOQ
q8c7HOE/5WKYKede5f3Z0lEknXxeF8Dw74IFfZ+m9NCIe9689gi/5hpw4omZ/f5nVZkzmlxWxbbZ
oK0cR5ThdGECVKbOaG9pt53CuarAbCDa2wgp4je4qXuLq9aE8pu91JS2eeRmjYCDQjzUNJNYXseQ
otBnjss5Hc2znQ6q4CN6I2eSUgDblxnCPR78jNP/+2anHhLq7CuJ12HNsmyktrYz4ojKBtAQqG2U
yu4Zweo9yuI1bTi2fu/FcZ9dElnZ5GDDSKb0p7amIGloTp3atFsyQSTWlLKYRuJe66mtX+fFwlAW
QUJTZf98qKqPenjWzzQH2U8qQ33AbM+GUgPOrctvpm/gaB84jtgddK/eQvrXEr2OfOFG9doFP0pl
SpKEj1s70bmskAuENd13uWg0JYswwfKyArHcve2r8fS42h8R9QvHdBBBKZmTEo52pF16MCI/4tA1
CRF/QaogP3etXT5DJmFpm2kCJz289JOQJbbwSnsS9NLVrKntnz5YCQfDattFHcyz91O7mTG/aebh
BzAD7vyzADtsoJAhwEvdbUYJ/w/xE7ZaGWF/BP3iFAhVOuqx0p70JVGXk9JRk6gxPIGaVSmzuJbX
0V+g9iJRwRz+KEiBdmnJr1NjJg7/RZQqZGoxJ0FUtqSgtfciHo2NqlKY1ZXc86p6tnvMIe3PN0eW
sWcYDa+98eT0RSoQ5vIvSNPviHDb/e9TyIgM+DU+AKhinKRcQvpIqRR6Nyzy0n13h2BnoDE9P0o9
cQjqeeO+6Louy8RsAW41mNgFDXhI7qdnUcmSJasVidvNhH8x1hUAE1cr9hvtqC4BLlFVH3v8OAKI
phMcZTXdWC6KdKGxRUGlkyQOqQn9KXO2/Pd4aaYF3HNaNtzZk/NEbFyNQW2G5m48/p72EYJNTxLN
PCdonNKHs9CxHfwDJZMzC7Xdydc+V36SJvl9RHh/uAD9SSthBVnqmVKBxSgs1i3J8v3UlDLVYenG
Aiv3Q2XFhTcZbjUg01WP9wEQUTwgCAYJ2Bx94IrCqnH9/kxrktg4WfCizN7PeQKjTvnkqa+AlZAw
4wgWPadhMnIWsvIKlBc5kXM5P5ELJv02uHWHodLJF9NVJ+pqVx7y718QakVem6bVtTa6EjfRonsN
WErcWry/TKxG1l7YmYVejjGNkZkbidCwb/JZtjmErp58wc2xiksBI1l4McQdJqHVppu6NVVVQYt2
nXpKC1l2cNlzZYhGrqLicmnE5H9TmMJFMD6C34P2a/olKmMeYFp2To67SnGFbKplZHSzqcTzGRRB
7E+/wFLw53h4DX1qeZcZUoDMCGizXaTqxz3heMH2GsCyNretuy3HAPbpUXksnVx2yETsS5tDv4S8
C8AOX8WtFPQrwoNH9neBatNRm53kAm17Wq42RVbsCDXklT8NwEpgtrNKK315chJs81UZP4W3N/Ru
bvj/59xf4EBOzgZBJHU/+RqJt480tOp6XDVIzo9WQwUW1qt/U9n+87+iU6wxFrZGpgNJracIHM2r
xR6pFXrxmgy7iTtnWjj5SOcZN3bjrLBwsh3zgq3tv6VLzwoRbJCFr8wn7YP13uWs/F/mN+jfv2ck
6LdRzvwX2PXvGgiSTn4em5l1NKrOqZH16AULIdCYnxyaJx9YJ7jQXC15fUSHrlkTT0uVKPpyiJoJ
SmlHTMFrExQ6CvrzCONqz8pkQCIF1sMm+QCcQjvc3orpd5io/hFzWfIPa5HN2WvA4nEgoPpZ04o9
0GGzqreITnNqHhvzy5b+L/Jxcyn/+ifUY/hZqa7RDs2izZWaGCOTZDklAb9vv5EhmQQrgpfCOQVX
R09qpQJ0tn9loZ9k4LfTDpiqOkGpuHB1OxfAgFZkPPBKQRBH9I5uM3IXhqkpiOM0J/VSiDy5PcXH
yIHsux1Llz/BiFu/6zm9qltgKkIR14qHP+NKQizK9ThuiCDAcICPqwFzFV4kqN4ujFdr9p2Tg7kv
ssujsxQVqPYTKbin1nRFdUZ1x/HA+/VPSR211AA7e/r6JXIhglMC/V49eXCMkbl0TALsB7zP4Zlk
7xRib0qwAHL3rhL09qi37zjiLsHEW5wglNyduSRCqFuSb5u/Mscb0K2uVlEzyrZj6kisCp7D7zfk
Hc4F0kTyyalE97J8SgfjaPtehWMz7JZV42PE3r0D1kSwefF4wq3sP+QdJM1yHgX6muT6qrrWeyXB
Z7fHNvmtiXhyy4uVGEPZ5lfYu9IPuQPpPA+KWW3HCdaipFfAltrdUg65gMn4+mlMIXX4tCgW3IWH
K2jVUD9zMlo0vDsyF2QzrGQa4gl23jvffZuk8S8GvegoQ80jHxlwqJp+8dbwNzeLV075SYXVpzOO
cBT62MRM08ZMa8es2hhftak1GzWcqX5BMYFvCTo5C1hHCgjzqD3AAtbEWzhHmx3QLTR1mqYYamfE
lrQt0YXE6a12Q0Gb5aSI7DpdVtpNZUFGNz9FtNWbWbHxyj87WrLJGGLGvkbE4/+KJdV/InR23btw
JeHkYw/XlRJidT+0v2gcp2qLdFnu5ZnwSL0ZN/cyksqIotEt6dHllvShsyroXY0CEIa1MjELvkli
oCJJcUeyONJ4H1JfW4nXiseorlellrzbh6b4vuXRV71sUs9W/kjswrUYdsK5cO6LFmHUZ9uhSdvb
jMdKcd9Qxh9kJIgxcclFpcX5MmPX83TgFwXMwTWc9yRi03PldZUYIgdABXw+MTMhOKVPf5vAg1Hj
MsJ3u46GV0PZ+RXDV0x7OicJ7WIiNHT+kRbimB05xfaL+wLSs3Z2B9hhmJ6nHzKrpTts7CuF7Wuf
dw6vSICaB3BpzaCu+z5sVjI6looCo/lfOxGoK7qRvRCIbnLIDKHR2w1rWkZD/wz8gcMRn/q7xN1Q
Um5thk4vIg+x+bIdsEQEVKt9jdY2ME7zdaJviSh1KKZic1ASYao7lwYqcgK9mjpve/IIn7FO5dPX
5swGL9qoXhjPjdQ1XF5j51GbtjMIWKQ5PMe4So8LCIgC+fVwtWTJFO0QQ0LwNWSGAE4TRqGJ7ct5
zliDWsAs6bT25eroBc8TqmH2Klc0uAUXSKSpCOHINShO+v0/EitFfWYVF0NAAluyhttMeSCnKr+z
cP6oo8CFE00KPajlbhnd/eSK7Mo0sqT0ElX2QBrkJwNU4p4xd99VBY6FGe5VQTMDYHDAJbtB/N+p
jhAGKcoJob/5+dBi3DVcONc7qxJrjIRrQ4EQr3AiwwJ4Yn7cU4YJd6SKZ6zKHGDkqCY/7d6rlPES
2JS2c0dAAo5xutT0FEPBqUnK+ahviPWMCSf8ALapWOJcbZXI1NXUmIux9D55bG33d3jFiaf/bjHr
4B00/pnGE0YtWd5LQuZOp5T2WE1e69xf/1NxB7+BiB+1J6VTCFJIMVXZm0/QH2nfeu/mqWhJlVpx
+9WUVRDP4+55G7urihgqt/gLDVI4thiN8gn/IflXzDZKm6UJhqa4P0TlC3Yi7WcWc81j0Vaas+Bp
NCT+LKqGRM3HL6M7YWaJHTA87fieryfHYpiVRiqxkRBwgmsCfFuo3zEWiO+tyRAq0gp4OMJz85oL
zb+zus15+kV07aANdr8Fw/fY43y5xQFCvF95s8nLYamimuf4gJJV2p0Ys6coD4bALF5xzJ96cPVQ
48+UtrBS2Xe28sP73cO/7k5Y7/TXP6rCDVF140bL07T/3pTgizE9SxYarw/wpFE/9byy5+iHDcZN
qgSYZqrmZFQ4P6TJd8OW361mZdXlwEq7/UWS1RstDL4sk9HuvinaN9CUckb2xcL0PRDJHDA8BnhZ
46BkVmaUfWySBx/wcU0H2EhqELppDsx8Ek9B5Ds8zLrkGoRyoJr2ExdoDjGn6BctwWwLJ9nsHogH
dZGjFqWJS6/rmrNUYW6UZtf/jEJDbcskyHYGhaQcTHSv6Mc6EvZMxyOuVNfSjhdO7XsGR6zH0yua
m6Lc7lAyNGpsw3WYL+O0F5xI8CCDWUgJHqMLrS48JLxxIfzjAbrhl3HUwsWjIXDZHRaJ93oZ1UCx
IWEBt+Vbg/1rjn6REAcy/sXjHfiMwcApF/MK6JTPqTAhRwB+VP10xjiySZYItmZmct+m/GaUxrYu
uKyM5ri0fqKpZIvmDPTQqB3vPIVWDncDnQqgbBvVhBrzl5Kae7kxchkRWV/bxxyRR04tadBJDKHX
70m0Qx400+ZcMp6nRGgLn/NhsH2HXvlvR9Dr49NwpIetcNKvPhMvv+QNgq/Y5I8XLMPvENfc4Prl
obpuQwAMlWRQ8BfkQvG8Z7OqF77M7uIsDH/bhTdCZvPw14EvSQu7Po0s9UiYI2roPeSKVIfc88Dc
1RklTD2ZWDoQ9//IGA/D2jmsyyUKlwuYmYCL6vf3Z7IpLdlizW2RR5cD0lso+InpeXfWPkWnZJqS
yYXTGFsJCjLLGeeFXL7Uo+OSHd7BObKeBaE3kKif2codEIuZEz+XId7P9ItC6rNuZbxKtE+QHUJa
XMeg27ez5o/gw6bT6ZLnZaDHImfZ+9tfuQZX4CS/N1scN7vlhPM7WA7Px12OUbfduj0bgW3yivsY
optzDlBAaupLRriFaVhjGfPoC45+nxv/C+XEq21zGlifuMj+Hw6EV+0uBJLuwSRITikr31jYWzDd
DEVP6nB8+aYuJySmqoFHF+lM2JGLGIgK7TG5LHDI+4yvLda4X30cs+GrQ18zG4MyfymxaOi8q7pJ
n6YCZdAzgfrcSfKQIDbd0sBZGAs6V3Xop3l9AO7oU7vVrefAknsfkwk9tly8SUbV9qROKbtgolfC
HE44vvSFRXT5BMCr6CfWoc35nJzIkP0iUggPWitbF0yKkDreorkzy8eKY1JCBJ2dUTYMbpRJ09YP
DHfprnQArAW+EtEn5IDUQsPMd6EEYRFuyp+Gjolllfjt3mWH/1uhScniZAnstJY3QORkloRzf1Ea
g9gkYAX2lfD7VhLNniIsjEo7uN+NVElXaRpPfrs5r3u5ZIqW2PKpLKxnBvGYAJDi4W5Sf+0sAmZH
RK1C52QtCic1vALKiI1DvOxKxCSI3tdcrMZJ5dgAAvvxO4w9urze9KoM4CXuXtz/kbLgZoxlUstc
WvW+404zHKcdurmKOywipEHEu/AiBbZFUGF2+ShAy7Y2OehGLmrc8iAD9FyuXytWziXgQV+vcA6C
icchaP+Mx5Lfj4SCaj/QJxmZbiyvMKGbLW8AXypBY/le87zrUNVDcVogzvG6GAsFfVNH+a6zGKFy
kAAflABXsZl46ZPFGctk7e+TLvr1rwavJh2rqGgk393AYMZ+IlX3FzLbSHfuzx7ulg6Hs1zN9yTR
iJt7+ghEgHWtZWy93RzzCYY5FSV5oS1+SS3k6V1iGNPG8ZGzx84SkViBNgaQuV57UhrEY45yQcf/
5742KB3XgOKeZ0pIpxOt8YmAmTvu4wRvWMRLhNi/cMDKpvLFL92iPNdK+wKOyZ9lPp5v078Xj1xu
2TWAF4wjGr+ucME4GB/eLhn1tC8LZ1C73K3EVKuRN9szABAz2Qp1Y4LxmL4gc/Wcb+XliWV1x0JK
an/0In+unz8OHUzODCTN50Y08Glsc+EqDEsoic8zf4ypVGFeM/Diy5YUNijAlNUzwqh+HqcmAKST
sDKdVBg5TJiIOw78DCvwrw2ifcQxZOLMd4jgQXYrBtK4lLeLXIt9DfZ+H6B+Cg4B/W/a7TDV3g/B
JBHUUrTokIosM49ENkrH99gOCK6cj8PGK++pTSZ9+bpHjkWUWN7SIVGa/QkBzMGgrKnk1utxQN+V
TKAdDROEgWimjJC9Mys3JwYzy3eA/17M5kDLZKkk3X4uQaKPYCwS11gHIQvWVci2WyqBj2K3mRZx
ZMUrxnA0jVZTzqEjy0+hK2JWY/3dGkAKEROKc0FCxz0rAS2lDQe3mRHsMqX4rkwwVRtdOdVVyx1+
jfRLRiKCb0yganhUR7zwM+uBnNTdI3yJ+G/WQc/pUewsaXm3U8dgdIqcF2PkZjQF2/Onb/J71MmQ
fKazWXKfn5oJN8477sqGcG6PjzvTt4SrYymV713WvNPHCokEHCCeGKorlFPpJ/OqP0i4zkK5Z1mf
1x+OHK7MROQvs5xB7A1XLRog+utzNBA9yRYflHWel4wAMM2tgk/luSIi7ekuXOCSf7lYwGzLcUZZ
WxHdUSBrQNOre57LX/LT3NvQghxiJyZYBs8zJbAkLG65Oh975RWTYdrtfEn+hCQ6uxpin9W/7tMR
ouQl3JXswYYik/a010lAzUraK9GA68yiv4h292VvTF5a5G+zUAJFBaSlWpM/6iRxGjxDIyi3o1ar
DtbegAO60R7/XxlXjYgbRI3oaHFIb4hCRg6+LehyzXSTmky2UucrZjI/Ww8eyyme6Z2h9O1w4xHy
9122B1JLfTP5YqhyeMPmYzqEnEJCS4wySGTTaMGShQ09bs8G+4O4IZT61DkvVMl5IYBsOTwGzQ3x
ft4sMcVQ5pLGuztyMf/4Ht97gRyBax+zKQPA70FA4ygQCFnHGz2m47LsvMgbQW5kX0IAL3QmZY8d
v4r9fCYqXJ+hg69u6vKAfTga86nREL7H+yfepesnf1od+JvZyY10O/bKiq/ZsbibZ28EX/gVhKIU
dS9u99JQ7B8MyZF8k3xI8PuSSASkbWZQcRsc3RA76LDxOkGz2FIjbNKpsvz953Ky4c2zwZPKdKFS
a3xORxUXwbWfjzPFEtz45oK3Bauw1b/jKdMVsyCg2fuIktHfp98vmSbi5Y6w4+0EpOcCZCFLt0of
GO6HGlUoDBPuq4ybvOCoR0zvETUYe52JIjuJb9bjFNSEg0xooALO841hYpQaoD+Hd0fdLUYf90VR
AQnigwS4JTcn8g6teKvvRJmlN2bDLNBhnrvHtaAComlW3LLMz90/yMwnRnMcZhbFeyHkOD9e5J1P
6YnEKPioIGjGZBL9BLGPHmuxufUfCIqqajINdiz3AnxJlH0Kzxv4DGsYFDcyz+WbHwqZOcn5NvWj
OSI6N1+J698JfY/BQ3ZgL7/ro6TGI0VILhv6FLd/FR6oLGuAafLim8vjS+lhwKv1NMY1GbQ6UBX4
vCVwhtLt3UY+fG2pXS/eOPA50GDtRF9uZysVmmufis6ZviwfLtVG55wy6aMaR7eHwxJ1lH11tRTL
7lUNBQ40u3u+2HoG3eNgKtzNDd3bMgbXM42g+ODqMaXyyazD13hR9bUHQLU7yJj0jniM6DJa6Zii
zBNuk8JxzO+BHi6NuoQhqrx8tbFe3Bsu6LaUBkzABcWoBrJ3VmCe/ur/TS5FdGmP6NjBIU+7T2/T
h6LGE7kQ9wcntDuydMIzvUegjDTPuQ8fu+xUS3SlQmI5SG0ZONAQ7v/lciNGI0I+xE8lHJOCSCyK
zS/7haHwDoM9zx6FNJxAMud+IE1846wGUgTGqYsPS9Iy6Wqc4U967qIDi+7fZBTw+eUxcYhjuPqb
YsEWCKa8RZ/4gVEwghR6M8DoKnRYM8h+lQVGHhSa6PczPYGQ2eEdDh7pbfpIPJnfrh9rrkAWbez5
w7Blbiw9zVKUkCzIQ+KhXrg85uxiomhgbFsSQMZNZqsF+R+/IRzIs4zjAHue0etKpPvIURWDdioF
WMO+s7yJwSz5xldIwE3ncqWyGGtJ9KHbwFn+DKy3P8lEm5he8KwMEFdqiTe/h7MZBwZhAxMTTM87
7ImkgtEWUjlg7cozW6kQTc/NCqWPOnnVgk4UwCebANjrcDwIARfi55xSxcO631FjOa4takrldwnJ
ZiTRC5m4kbLyTqlHmkj7zRYGHqUNTg1fts87nnJmGHpuXy/jrFGeqK0Ax83vu4DuKQd9aXcwWJix
qm1OVxulh8wL/QAKzDzyP2J9ifxsn9VFGsTYZzl6S3q88ZEjdVO2Uu/0s87khLDKNLT8FZW6a4Zk
/898epFOBwsyWNWdUwx/l8xQRiJEquZ+OPiw6SEbPi2SNeSQ7f7KS+ZXkHbFpo3VU/33xNrF7xlB
YWDXiLUBmTYre5aApXEPt+zKVOAzKNAhVskcxKumK4xtsv+6SBGu6M/M8CXjWnmz0Pq1Rq1BQACY
C/v+xYLErDOdxHACTcuavZTFwvyT//YhahNOve0hcHxEygvNSrYg8q+HlA9PayZBm6iM8qiquZQY
dNMxsF+5dpiml86vrhFrNPeSp2jtL3tLJ/YZwCfRnSe2J185XS3RbkqMmwfmKy7td4j0v2kf3oWp
dHNX/jAAJUV384CJ9SIyE4trlUs9hGgVGqvidSonDQx4znw540AUPH78UYvPu0mxj3+Mqcwrf9L5
/WV7maCT09j+AWIQ1WIDXBH84bKA1Tb1gytRuLZVvOCxUv44rWpiriuH7nNEfQlevBdQ+a80XT3Y
ycQnBVJJbDqigJODcbCm2m0XMuNVdnYc/Z46BlPXuxtWKCkf6bzYUVtM8bLvmx+l7BNc584AaHy3
4thD2ktwh9weNiE1T3PXFiq4CwEOX6zOVQKsmvzcwf0WdJtyRZvfGSnyTCjBeTHQ8i0yvn2ZjEok
6+WCkg+WSq7PF9wE+jlTZlR1vhPaTLmSpnHTeLbnvEULMEEDnIpyYCQWMH+nQhZHfOVL6wpeh0UT
+n9AzGmJ6V74VD7WdTktHfv6AZ52ZrNZav6U3qAEFe7oLPWUlOoKbU9m2yA/sPa7fB/qamSTxOO+
7D9vRGnMNG+U5R5zlHKnQnAAQ/53hl4ai2QaO9vZPZwJT+FVjgHNKGoHmI7c4hQlbagqsVC7D4fQ
e7TpZa2Bmn7NNH4V814fvG+Z6Dr7ImVrCVXRbVLK4/0uoLFbGgZukL2jC7TVLJRHM9Y1U4JQzo/u
N4pQzSGGWSIISfkwp4PqzLdzmZSgwCN/aRSi41yjhM1C0iYkQ1BR0gfkP2P/GDB/Jkl/CZrV5mk0
HIv2UQYtGYU7AyHk/Jacp6R02imAvww8mxUVWpugTGZhgy1Et4bzoHN73b8umgRm4YDN41VzLY43
vrbS64icnLkq4q9SFz9Rsxl9LEIeztTM9vXDNksUo/b6kuZ9vwI+H4HnQE2JV85a7rsOKb4jFFvF
PDqKEWQGnjvPz2j4zUjTk2gMCqVf5m7I2MDzjx6e4u/zOdGVGOwtbPp9fuEyaQn7AGlbTd6InvV+
Ipz2wH+Q9ZFs4SQWeTgs084sPtiV+3Sb9RrCuwqfy+Vpc9EQ1cYmTTMiV4b94fNHuO5g3zOb8FJi
+iACQ7y5dtFDWlslDV1pe6GG9xep++SpTBEHPIYChn0DgOH7gQ9+yG7bc/FNVPmIshB2H/r/VyWy
Tzl455JIOq7DaIgW84dt0jVK/uJDrHRqWwfPEZFhXRa7pUh+BMqm7Q2AzIqs5oBHhEr+ZxjwSkoi
qf7IcA9+f+4ja4mvlWz4ZibzRGGj1yqli5cSVnFwbKMYlf0IOTcCcygc9cx67C7F8dAJjn+1JxyQ
XCqh7SSXjDOThvWthUh2auy5Ih/fTeSsPIE0ryhdn+4Kiz/6Spz7J2v5hxsJnC/0Ov3N8VhNmvTm
NmfinoVAimtwNDMqiMRxu49nJCxB2f4xJIz3rvZtyJ0k+wCJadGiVACr3E9UmDcXucmtT2+kUO79
YszhdyrqNOEGVdlfxzovUlZNa/brT9K27E141Ycu/+E8jp62MCLEDPmDsvfdGZ6nN+QTbaP+c4Gb
aLV5zkHu/EPIS47z1PaXNpigL4mI5jwrAcrQ5WIboXmNBTbUtJn7DccYOfMrnqRe8rnp+OC9vB/f
V2Vh/IBvetKJkbk4f1mdhlOOs4bD6VYd9HX/CYxpPPsY0vQUBdPW3peqVmRddoNnM/4BibQdcGJt
Zf+nAF2ooDZgT2vhmdgtV0vflhHw9lZq4ysQVCObBG923L3vhmw+cdHk/yVUeOQ50bCo2qymxN1d
rmgzMYTLe0hVIQ/yCSwY4BV4l1YiUoVW3hA7mF0cV1OtZMHx2p5TRj6S8RCBBYqoSg/R90mFqERq
hz6RZXeVLCBQhHQUlJ/j/tvuCtO699fp93KU0Ge5JUymigQqxZ1xNRrxOaFA9qEmE5W1FR1RGFXC
RpzwIZe/6zclOXF+EBZbHL4RV2BA/kVJxP5scp6HIlMt5gUG3PfWKISNPjOosZWmt3AdZM9e9z7c
q1k162eQquFJKNfAT66VD9BJPt4LmXYGbpSw4Dv22kOEPU4J4fdBXd+jaq7CdoXSGo1TgDG0ASA3
A2b18mdi1BefAycBqaeNDLJzoJ/YEfo3XTGZbUcd1dZvPgOI7yaC5es+yj3o9Ap8C8ajsbmL+yM9
QwA6QwuKIBclTfn84TaQGoECozZE2V0AKWgesRimO4Ir4I2i6BeuIz2mwBvN6S6XhAkOb3yeiHJV
LrLbyud7YfDc9iQwnhdUt92IQzfd2UiHS+wP+dWThfufolOsHfrDs4s6JE3InsX0IQMSyAnKaK2e
PwouzRpCUFDDA1UsMX4jotgxHQml2DTQ2STn0IhWz/nerRSS8KyeyIaTnu0StspoYDzhidh8wqYO
De85YMDDGG+KE4OBttkouwBEMT7DD1kb2b2hY8FeGMS0M2GpyE2onRQRphhQLv26m2OQLaD2i1o2
ETm3od56OEiednkKlfgHcTTb0iuMYi0SW3d3Q5UvfS7Li+IkieWeycSTlURR1ihDSc/yRQp/BkCb
aC4MqtHJ8Ss9+tJNAyZooPU55WB0OBfcekUCIX8arjz3AWiNUET4oSL7Rq+VU1wK2PFWjpjDARIV
4nO3dxSpyy7CqYkyyNuEnSx4Kk8GEaTgvqkcG6nHa0PmNOkptEoc44b8oZdAYaAe7uTm+krVuV8m
KAwQdg2dQxqPwF/2qB4cGzQqjaDltq9GwGAgEgQy2l3SQQ9u6/0O4jfc0m9fh3XT5KnoKboTtQTE
+iGZPni5dhm24V8s6BpYKIMbaprlHx608eEYrQCWkNRm7AU03hUnk/aAv7rfLevVdGI39beVZP1V
OSu5MJW85ZQgcIkBzkpwQjnwNW7foNVXHRisn1UpYXOwIyUFj/0syusFQ1lUdjJTQBb38bwVnCYh
dyDN1yrEXgCZUedBD+SWY7CBCnyuPQrgfN3jPaAZ03ruQBqgCL0zZqFu6+ovU5w9pplvkLJmfmMc
FwyFfWERhi3n/velKBetrg/mJ4tT2L9Hsgi8WF0zn0nMA+jXsgPyf7J/t0l+KP6NyFLjZ/CoLksm
YGHayc7MkozRkW3CNYT2iEBEvkobcWkT9OL9YBiCwyl0sTJ+kydwNkJy3sfHnagYEjtL2zN943gq
r89UeobYUEyZn275Pi4vAQOQRl/a0RDPzNAK3Wk6c5gLdnqQbMh2Rywu5z1UjKf68cZRx/ofxFbL
pKkh3bVJUCXLEWyM9wnWeI4EV0EHghAcRU84hJyv1OaTx1HEbedap7lqnfiAFz7h3L1dkN+raQim
tEznOYkpxtqmeYpmdnwvwuQzyxFUJEd62l7EIbzMsFxgS3W+aVmLz5+/rQfj/sCB9PMjzyrQdzaC
ZNJYUsbYOC+ikKMoI2kQdEF3DNGiPJ5tPg8ZaLwrvMqYak3u+U7JWdlP7LqxbkNe2ZEHPnP53zty
/jDjzeGmWex1Fd++E8SEyjWv4Du+3Nr5Bz9CTIFjFT9IhTbg4pc8KsDtzzf9p4SNU8cd38jPSRQg
n5JsAGfRKD4otLx7IE4Ptx30JqHgm7begE+RDbsE6q0gLXsyApz6hl08CYpZWM54/68baMdcGydD
EJZbxSLNYQDVBNQDowui9hSD5FUVnw+sKRIYhQG4l5vvS8IySXY5pkfa4Nylg7Xvv7t+lNRK5Lkv
MPfrkFGoNT3tWqojSbfq0KJ0v0LQv/F8QpDJtxITJ4jxgnuEt3wIXKcuGx9bIJclCZ1rn7iDoDHz
xWnimr6cpbIQgkjCJwKWcu4KHnUkT1uZJiCK8oBcIwWTaDO5VV5gdydqsASJ05YWM7YCcntPnhpY
msbf2JavflBKLLCv61R5QHoWhcaBRgYKJUhX/TR7ZDTthk+MXNmWcPirksRWBsNxN4OpIc8CQUQX
2+/t5K0jVdQ9oMWdf8BaDXJ1BO9BsgTmykVnb4kWJp3AQAdNjYwyRsEI/LzlkERVfFvB9EWkQWFw
77Nq/HEUK2g2XPd1JSrHG3SDmWeDtw1amnue8sx+l8FfklpTIPzEOzA4vLLE4/dCSBYSOZA0fbnT
m8FgfZ8oA2x0Eg9yeZGxihgV/LgaLnTEbAsxRSE/rrzR6jt+yW8F+OwyGIni6Otah96QMfB92vJE
uci3csmYTPYg0HTLz066BqchmAO0P/OkIpA8GcLTZmBXN53FRFjRS3pyDxwOGJuD0GtPo3cal3Yw
7U2qzuwg/YioGZpaTQ2ZpZpnU0tRS3baA06wgo+thtzZteD0SiALgrFdgXlvWdnLjs8ifhTwGqKE
xZO8n0tMsWFKBvyoI3Ai3klOnF19QjFlVWxpA2j/532fqUBB0GeikmVWbzG7WQvDR3QIF9vmLdJ2
mx9t5A/1F4gdpXaAypJ/RbIAkU9npJsz9BpRY2sLSv4fHOcHihy/N3UZNR8cCplJI4Rx8eO7qqsF
p2P3dJNjS+8n6FB79rHYH+lAGthPglXFIX4R4+PxPzCVn8pyXQ8n5WJlCkmaWPh7SQuHbcniMrP6
l6Tn2LUTn2gwWaMQFgNN4D3FwTU5z6M9zvV7u3qwSZLM/g7FD8czJkQwWAuwKQ+MDul5qh+ywrgQ
WEVJld9doIXPavfBvB7VZ0895YC0FQoJ12RahecGklt1QF634mvjNBfwyk7ut8iA0lecps3qR+ZH
r+yuz0ptSBE5hfttlULEEXMKCpaEx1vETrQaYbWe2N5l1YMH1GUAAfdRpZ8NzfKwPh+z09879DkK
gfZCahgSrBPDefQuaDZfNQ7zvlX5iLnJRrBfQ080OEX5w5lB+7P8VT71Pqgja+yURwHqUAIliqPC
w41rXzF/zriHVf9BxDsfylr9rtObGH+kvwJzuHpzCRCgMf+5MT3FtVxIdoE5ROUS66KWNEVlmTzt
QVBAGH+w0R0jiSMdZhTdoKIxnoFJ3PwS3ea+SmCGy9FfZgEKVA2o9iN1itgmNsoJJxMmWkTF1Art
CKv2sP/NMqW7GtW3QaawTSZGMLeTAhxpTS71aY0xtS2XGLTa4SnpCocd8KTzoEOJKg/FjZ73W+us
n2JTUM0XyPo43ky3tq5u2eNp5ADuj+7LYQ9Pgh6YOqOWE161pOxoB0PhT6GLKA2g0NsBvCcL15xj
OxoOW2wXzGffJCUO6NNODAcjEJmOiZYlM8wttZgDf662mbMXDbTLbqhQdI1v78PgjGPgUivKB74B
xqYegHjNcLV+RxtqqdFhhF/TQCiNN49MRED8fkynmWmf7f+27c6rg5+jp4g2HEJNWwCIPtpNu/51
RPF65pnJqU30+tNGonlrmy3rVtSVqIIdzcEq0MY26AcBf6/2Vhths78KyNhaCnoszvuK4vlKX+nN
XKlNH3PqY3/3na6xfU3vQ0utTu3bobbm7VFgGfhF7xHnyD8FUyZavBCJAqYl2uG08WNM98su76+S
cRCTsPfIeJhAf7BXcrV02XdDxTnn+5YbGmRLasizmtdIQqvj1wDDXeFVzCEcOcNY4FV6ExDQ6Y7p
dZTrISfykaQaf4U0dKC6rLLzwgV3fESUCJf+xfxBHGDyoW/8rhOj8YsHdd21PfpB5/vdBphX3GXt
1bzTQL3vwxUdGo0K1Jlksxa3AaciPuay+xXJTonMVWXkyGLHcoBQeHL0fNcQs5WcU5bmyLZyLlrS
H2yuGvY9YiZa6UgCK146Ly1s6EV+pNNs5Qk9k+lQam824dFM5mmmJ9up/HAkM2JhOZx2YT+QO6O/
A0KIsEi8+0Ti6ilQMXUJTZ8oRSKZnr58OMhV/IkywqCcw5J6n18Q+I9GWlDztd5i5D2/7HMOan+v
gOPbgdEhHOIlZZxOS7nYoixuepTkAihQhxBCQZ81TV2T6+xc4QkXdpRFgh2wpn+4f6jPvZ3eqHeo
3JiaXetvQHhUV6NWkfSxml1L9FX5DiRV0AJ8KEd/fPpAyJSbC7ciOW2MMwrvRTOkO/lfttBiP5jV
2W73rO6nqNtdVExeROZ1CkHSmp3hZoYeMFbxwg1HsjsHoHW5/cddlKtcioPgLSkVnhoCyw5ZmENc
+322ax1vq2sPLWzMgH8ObwyDOhin7vg044SVnwPvssW1tdeDNhWWG2+6juxRTahQ3f+dKuDA8jjt
HVBlwgbVPOfL454nssygVcI/6UT9jC6jm1ifJds5mj0kgR8dAnl9RFILf5AI2/qpSoxaEkQGKQBH
g2YnLcsnf2TRGIUudZbcrNPiWwHkx2YwSIUkWWRRgLGnCWnHFHB3Yzd9isdhUJJU0ix7Kg7JxBhZ
dPuO6rJ60VCP5ADpzfaloiilwk013QHD8tE9P7BEOHLi4syureE2y6P1XHHZblMFjGdbd/Szf8Tk
pP9mzcfQGpvyzxu8bzEJ0zHvwdyOnGbWVD8nl0RFdSK8g8XvAVUnrEY8ic+jhiLHgSrTyPFHdvd0
5MLSgffOBq/LXv0xPmUIM+EGJVyihcO8HnzxHcFpKF5cX8j2VvAESKRSnrOfamGgQlsT1uWCS2iN
sR/MqTh+NzJ8d66KpUstFild0StvRysDbu36fhVslWcaoSuyUJzTGou4m8jOVhh6R6qVPBHqd4kb
e28ECDJnRsRihZZC/PwyEPR7shECsfQOgyzlpS+rbJ0U1J8tOm60kg0VnbN8f82LWEwvPhUAxCRO
Lpabkr9iZe+uP2X0z7meMMCHIVricNfFIZmt7rLEJsBeaQOq5/avUDYkv6Wt4NVRXhAaTMaD6USZ
3ppLb51xsZMQ2B2SG5A9WuoH/Wberv2EUXJwxy9+SubHAvRrHq1vvY+e82AgrbY3d+3neqLmpyOB
M++NURJW/Nlq4AI8CnjIX7IWmOu7swCebKg+77RSlu1AVGQ243TpZrw/oKjE65zf/nELR/lWbuJD
SAVPpgx/h/WyAdmltfe5EeOw79B2gYeBYz57ZwWRU+Hjry8l29sRQufQE85R+ql0Hg0UV1m4//xv
soxXq+/RDB4R3UX3z/CmRZ+KiuozPmPLgLQdr6zc7vRSPUR824o3EkKx48SG6dC7glWxysF/Il4V
/i4DpAAfs6PP3HF6o21/rHFFC9tr0NzGiQF+lZGbLQJ52pwy6niHaERBZatrv94GPfX7lga+4MJT
221B0MdG21ZPB1me5ca3WvwnTV2y+s/34PlVE3c92hb4IWx7p0FZNfk9iHhMuHr8PhFw4Ukxsv9u
5TEQDyQeonwt2M35gTE9fasyXqv/On6gz3tS+Q7SicNoY/AsRHv56kvLmUjF8DHEiwK+5rsyN7sQ
YyTqTm/XeF+Qgqwzjhql4fkB0l1c/83fekelG6wMA02FsPlpSqsBH5ay9VddhkOPV8vuILJzV2nd
HauOl1toIth4qgL2lrTnr111Ovno7JaaWqkLydVdN/BLOS/5O1B8foqejU1oR42v9vjG/jlfwFbQ
Rq9vtfmB4QE3eLs1T5W4xZGWITP/hFDBPG7V1+aC8RBAXI82tsZ4E8dtYOBCj+Viv0SNG+qsiojP
hWHx0ER7RbNB215iGRP7jQ+X2RhQErTzgVhLdubGVBCSgqM+NqXvo99DaKKqczDaZN+X1dRgxT90
r10dE5vg+TqJsVNr4d1fzQakVERhDFQCXyIbmkT8HLAzAGM1iekLKyF3rvklnxbmN3r3EaDt4yT4
oVnYIxDcIa+b+unacU8yINsd2RORFHxP15LR7xnNkJPMZeJF0pkMrWjSdM5kZPm6eP57IP3sRhyO
X87ITK7GqIGEP3EAAWLCJ12N9SxEmVFY185Djv9s6PROYIyjHOlZYO+ptAK+z39pqTjnbfC2r17b
3/nyS+7nLohdu7IR70XQBurjO7ya7wRLl+JD98xJhSDoKSiHoxESujSYeKMa2DBAHnXDWxttOUH2
htjCdMz4Av/3qBrisQgV23HMChrYgVqjeNt+mBlbU36LYgZGiWkeBCoeI0r7QSizvljg7dzTCnMR
sFKKzQqgU8lcDkZMqIZZBSUgOTnTZgWCGm3R/z4C37HO//Ss6JlyWQh5Qtq3g5arSRJAIixfucQ+
8jKaxQOyvI1MzbJ3p1gaICxXWNoBYZz/H5jWQrmkDsObxBpqjFDmvBdVr+yFaJHuaNoUstmwdM8R
c4m89Vo4ufDYG1begsD9rXCsSN6cplI/b+CpPd5aUjJUhF0y4B+n7n5gMspaj1odq5uFY5VYeXrO
QC1F3GPcHb71OwLvBa7B5HVK/R1PJWOzUlDL0QTGp5/sqGZpY5qsDvpHloF74wOk87XX6YLDxdbP
HDYwWD0U5uYwT/MuvybgImJqUlX23kP6ZUJQRK/e9GfRxADRob23TQZHv3GZij/SIQan+Oad1erX
IRz8MMH8VkM9H5sJiJgsVlB8l3cjhBZxxWamkmXQwTD1xGeCVxi4Yw1aJtBZt5bkEtcFaxde+U88
ybGneLKv5t9J19wM8LtZSEsTotDyVNRT5YNus3Ci3QF4Xcnhokv4UJg6IKOuBCe9CytS53MCBF3E
tfwcJaqf6xLZw7AfLkrwvED0WOgm0kPwRxvmsvSJu5S9LID/k+oPEZqijk00hVm4EcTnrv2MfiP1
M70UaatkNhfVXBlygWoGNh/o3ubNp2xpg9IrdriCdkKc2t2fI5iPT2dH5/qlCdsw9VDgv9EgwpJs
LusHQupNye1yY7WSlOh43ZSu57Laja8goz5yjBf1m9S4gTZsxKfkYxYtovxYgpq73QFm5/YZ8Dqz
KuiDeZHdFCtAk9KKNTOAzwZJzhVlhSgTd0D+n12RLJ0WgLsx443QDgPRrm4X2DOB8xma6L6Q/E86
8qqXprCJzU1q3QLKHskGhCGvsipQqzDAYzwWGO20wGm39JBJKAgF9CVm6eB27AL40XXfa2LmOhYY
zUGh3yHhBArekopJUc7Jn7UOzRFOQfkYomzmFTbRZPKpwZMcMfnEjNrYVsqu0cnEAr5siBtULU4m
/muSfeg5j/YXack/5KPnrGFQBqSfHVUYEj10EcsPNibP82FrJq3Xho/CmWqbJxqGOw8odf+rvwps
pacnppWVIntXjJQEZKU8j7I1RbprCeoxnhZSgmLMYcOnGNvF8OiDKR3t/KouPRQepVBSOMIl8kCE
f/7nolHyoMvWFGYRJv1PaMz/0RdDQUsbxFzOqFmdRBl38kF+CE0D9JZr9hVTHXyH5EG41zpaVRXC
RJZa1X5xUsvK7/9NVIIeLaBJ7q3wwuyjd4dK9f5RSyr0XzOsvIY0qt9/jI9wMHKas/0MfAJJCmSN
mNBIG0RwIA2q+NLOsQ72j1Dor02Lx7p9SadtTURNv9TQ3nyqHT2tSUd0UkROM8vufOaNzRHv8+2J
njeqNVPvRdX3ee9OY2VeCOiv99pQ8GKo3imS89Eec0JrsmGqhzlDmmg/bQ6RqiIWe45ezpQMcp/d
Z9C+GbIq5nE3QPgioSvOCtHqUfGu72fopIHfR6elP1IF7Xm1Ab8szdLGvUuO+ZGrkx1cgeJCw+R1
Dk6s2i/Bb1vAvGTNHU3WjAfl7U6ciZmZbUp30DMvqXn+5IHNEcorCkdH/hJtfG9lpk0kVve4Q7P0
m0PeNRRJWHvgrOpYxbPxgscfB3qaggkZPhAF0JcY3P57g2s3nS+GyLDuotiJh6CSGsly9OMWwE5K
eSPkGssenX6jGfjwH3VnjAARX7viDoSMiqjL9DSuKBku3U0/KmPrVPAgptkOcqNnsof40WmvgJGT
QY6pl7N4ea9GfdonuBbJS44Z0Am7xpxlMSQZ7hvJWYmIMVbFZpFSCe2Jd3I5ZdnpFnk7dwlA1Ah+
M2i7lRN0NVt2Nk4AwGuo+vb3KfFl/59x/AFNTfrkdCf+K+2QQIs4BTztjvv/yGFTyIwkR3CQtZMW
LDpQxLRSNrAUFAQiRKZw6lOtqAAbRDv4HcAQ8vWaysaBZS2vVsiqwB7IQx7B9LW93RzJMVm/5Pg/
SnD3CvuMZQ8zAZyYB8Ij1kYjHIDBFQ73La7W4DGcLQpCZD1fMvoG9GoqYH7TwfXepEgouGreRJgh
S6hlnVkEPz3CP9s6a4w1UgXsC+adyXQaHusn1P7vQZysU2jJKURZN7CMd9F89lL+RJ3B1eI5y2Gt
YZRcnR8CDabQXm7bMlAi20GI1yjYZlMsnTC53OZK85p1CJ7zbyliW8q8vWSPhgO3PGuMBQMdLSmz
G0zsMgOfgjOXtxubT49FDemGCQ6vcsvPPJOcNVdrrwWj5tzwbK8L7Y/4RrsHagHiIobLr+CPFvJc
oAifPOFetJ7K/lsnBGArPRCKzSrSH1xuz4egOW4YD4FNzMNo18VXujT5admGBYLOyRLxmPvj/KPO
CTfbgjC6xbnvXe0JdUwopsPz/HooSXNalQtNf86/JZq1nANZHvG7AqykEB98QfCYLx1RZYESjVae
wWRwZJn+4Tfs0MkWCwKIwyanjHRGcT9wcosTXQ8aQpu6JSZ5AxsoGJZRSXUAvRI2IYS418BcoCLq
0EhmIqovprfa+04FfWSZ+MrQs66Tnl8elpKn5Zrwh8kpz8AmypzgzwtVxsLzBWcyq292oybrvCzb
K7jkb10sMKB9RWJu8c3l1XAY8V2rLTCh0PZKssBItQfFKMQIF00tHrN0BZnsT/+4RnF+kh004KIr
5Ja11oAAloOCOIWslxoxuKxKZI0Nne2xyZN0EwasYmDEko/OKiTwLKiZnvzlcvBlZu4mJNVEr0fo
WMS8UVPwibP4S6nkOgSv4id5K3V+0sbWjAe8e6FL/IzZP/crcPCrTHlRfzg3mbVftHWHGCLDHYh8
QAamxyPq+PfgdNFEGcrd1UCe7wPdtEHgoDMv6Dot0T64FKiJOVFAAhPCYwnwsWliV8RaCLVDM7CG
8jKB5PYz27a4y2aNFOHjLleYBcGDmQDgSah/HZ40UF4cUmzwptsgqJbLIhZSJKuCOz+EP1aXLX0H
QU1/7I+3OoG1iBKqRdMhJB3xjQg8wDVFwxXvkk1DvFPrmacnrHPRC8o7TgExeMywLBWqJkNpW07E
pq26r0QOPzPgu5XT8bKK5JiVE5/dc0TshJWNGOx+eDI2OzSwaxEtM8Qu5FNxvbEBs3EUkgd5NzV/
zYkX3FSLD3IJSv/6g4dQgGRoCLgY/4QCknJE27FNiTBTINxUIkYgJKAEd7ifGcq3JT9L63HuNr9r
NYnxboqGei48jl6GT0Fq7SgKO43PT6ZOorHaan6YhvTVxpxrEIA4wq56ul3piQe6mTY93JZpCLq9
KcOnF1h3VF+ZIRRLix6bmTJLUm/p+bhLa6ecBNdoqNdOg1YgXk9zGS46Lt6jRjkL8boozMZb09Dc
NKRCYkE4GxQsCbKZG+Le4oiBI2s+c/wXzRzfIUsn3EdclgHGNFE6iI1vRaY6Y7fIRk4OrlVso32X
JQf7z7G+0GR6jxM5ROpqyqiQ7Zh1HlUZswzbe/bZ/AcnEDUSKc/POI+QO4LNmACLSCk3L8YHiy0x
l+q965C9qhheq8abiuhdPN2yEqeqkTukNfwt7hsT+sT8dK+ObbBzcWFjT6jdNrq/DQI+3/ruCwSg
QFG+7SiHQHyYfT6RjkBnWefi20kdPP6HttnklW/Jr1aiG1o75IGayfYg4C5VMjuTi22bh/lKKZH6
LJH1GXQLNyw5SoLgre9AMG/Vol68q187A5J1r+TojrKXf47bPOTIpTkOPw8dyVd22AMFvIhKLeOM
mFdlbTB2ffSDXH56hCCsEw3Fyy7cHqATq1eWZi86jIitNYTnf0g7upaPnuEVuB9CGQLVvC3qS5bz
nMp3TfYK6s/xMAhEnS6mKlO3SK5D9ubhO+vQNAVWcv/qpLZ0RpkfelzfRZUHbEZ2COG31s8vptv3
2BNfSxNvBmwpVv3DXE8F1q7Um4MYUWX3roKAMGo5OytOFG6rOQC2VHFLoZRSXEHvnnw2RycN9JIr
MA4Sw3a2YjpkirjJ4/BAit8edgUWTf3GhTh1HUhZj0Gr7pnrgBqphGUaKSGiJPPdH1qeZZRZtYdW
ubouBPa9624m2Af8JPqrUBlvRn9LdmoZphSwAtzuGf+DaMQ5wca+MN/LvcJtJDv0w6aPZ5Spdz7Y
21QARkXiQWhxt9F6DqyHZrqwrWFfjpW8S/p+jfkI6Qv45rFV/B9CsSaJ+OZkQHzuBShtD1tNQz64
LNF5I5DBfRUrrdpWluhIxerFTf7x5f12xZ10zNSHdSNUmTlu7CVdC82Oo01Tka9sSEXExE+6MekD
x4H+SGglHE0rOqG4Fpu9jHRufARBgYp5b2ABI+m9UosABY5e8SDdaWwzV82XF+hxPdHTdP8niMrl
f2qs7kAGWUZR6F8QTbkholTIoiwN4OxhYcJDDe5IciH877dneuL0uaiyH42jLQ2lJR79pLBOVSqD
FwS1R30veiDThh400pcP6D5TC6k9R0YQemD6YUL3vLo3K1ONZ9j+Bi3FXZN05/MjKPUV0hwTliJn
TQKzO5DrMiavxhS52L27l8dCDgEGsjHZ0mftfwhhBZiHC9Pif+UM9IRZ87ZPi6l+7orxZUSgZAKR
8Kw+UEF+TY4sGbCUbYMi/3ubllKAW3E0lvsFdKFILDyNIfP1G1RRP9pCYw3KMPJfgNSIKBt1iiPO
4oMhAcaRltWtbtBeBxZd5HdFLrM88zf0xsGJiETl4XPAvFMZPFUWx6ef7bURx2r0IOclY/5zzq8g
YzSeWdv8RNU9Etbibf8qmH/xaHE7lqIfrh2XKlnMyBDSVo6zRqw9kDCeY8eeGQ/Z6HfPDQKPiokO
ow3TpGnUaFbWdB5pYW5irKtU6XgvdQNXD/Ks6yf/OboZALyBe9FG0c6dzI8xrdP5+jVXYUJHbPas
pP54ZhiSFRnLoJgZyHeYuh1KSuXDTiyktWKO1xqZWLC1Lx/PaaQx96F2rHCemdm7rV4KjfUQLvbV
20XcNuL4qsxEVtLLqBMkF8/tXkynzJxKAz1Gth+a0XSwDoBrHzUTLr84y9u1G3h3il4018aKRHHZ
sx9z6jnebROh+PVEDeNjLuG28XzVwKqwALLloJQU/XMxix/hj6Ib+UXLGX/9tBuel4r6McqEJFfz
GJ4y6/xiXXCNsJfZKsAvKA3SMa7DtPyC/pdFC1vH8UjU4uKur1PTiRtx3+7cxxg0Retef62a2l4x
VjmidTuFHVehqn0OBOsKvnZy4PZupwa6lyhsEMWhYskc1IhNksNXBjy9ECQ1yNAiYS2mAYVe3Lq+
GKykEVKJEOQzvLK0yoCfyoj9hO9/n3PqaFNetKQWUn8XHtZBbzLH+0R/SFHbelow2p/B8E6p5Xnu
YHD6XrpiAQ7/6BK8st6m/MAWT6QuCetcsm6PFMLn/H57cddBppd4dnv5fxeAxp7UJJLra6/ZCy0S
mpI3wYBuqQueckUR1qBHBXTNljjk03lx56zfk1BGW2pxpoXFbUuT6WJESGn9L5voFuiuIhb2ZqjN
BwMTjfXcpNnvIw4uXS90Mos0FguTSUnKzFESAc6AAY6cIEhiesiZyIeju8+8dprHTl40ugcRVprJ
XFW2gyR5FIE7VfHPloII1K4TAnt3fgzWOFb3HrGCriJIWfEXLOSeARPUJxZ5pasTTqMHen/iqjRQ
bIgFodkI5DLtHKCXZSrVMnozvGAgJaDYQ/xrSSD+beIJnIMeEDGNhQS35dkREBXHj0VumigpkPSt
bqe1RUkm+2DIZpFjXqVoQ+DiM2z4/DXhTes6UuY+lQnDftTyoHBOZ3jGf7egKvKCUVbdj9sAzZig
4xhyWtSeKSbmlcO0G5k9ZU1bB3pxL19hEJff9c+I1z4gCp3k2ZNqy7tdxm5LVVIfVt54G1APN52p
FWC74BkBDSgxjVohDuxFy7ZxDlj1L9kCM7gt4SeE1ekvaN8j4JGP6w9c0CKABawaGj4nm3lXFNUt
Wu8RdZ8j1DceXbSi0Fwb6l/+3W0ZQ2ylR8/VnINewKNlkEfEn8Gt+Be2R7zRJNdgBNtXWh4bZcvI
05TD2VCHd+ovhW6xczzZmOaTjIo//Jd8P50GSwI2hJQ5eKFmXTizm51Kw7zwe5OnZVEFK/03vOmK
/BwcqPowQOq7y2rIYvbEfZ1rbStdpOnbPW1X2CHEo4XBfbrHbkAQ68AjjfxjxdzLQ/YjiyMinLx/
UgF8ENKyX/AVp40cUZxXG4udMklTN6UyU+ICGaDD2IuejmvP9JoJHk/KMcEc22Z358KzSrKvGqd/
qvrFriPyxdefxc0qrfZ3tCT3AoOlaqm+5yhe7CWtURelg4PLXRKMJeMrxXDPYMjoBo4gZbugjx5e
3MpL8Iw85MihNq1YWgQJw4EpoKTYr9eWUJQl3zwmuKr+I0tBamwX1qtyK07SBb87jujeoziSZmV5
BT3TUrMmUmDD+dTKvPAPqrF/aXSuca3cvj/6AAASI632BOIAdZ2dnMHNT41K1x1DirihbNLC5Tb1
/MqVnTXXCZpPv0LVkAHWXvArO32aiB9VSXjVSqswVmGh7UxAfGIsTgzlVznb9EOoP30vJ4P2NlA7
dJz0QzP7P2cYyQVicGpYiCFLWrhl4pOaXw+LJBsS6rw2C1VFwu22gtiptpb6SnrJMjQjK1juUju3
SRzWkyF419ryxy51ZWl9CAU5vLdVxhgwls24ugdb9dUMij6HbC0GFzmGabT76YhMJBv0HnCPCiTP
3Yt4uKNEfgno3YpzJFb5JkITjfq2zlXOpQR6mWyKgFXjny6o/kb59sECgi6Y97fYRZ5m1SK0NwRD
z+P7vq8E5DaoD1jjcffTGwFkoSX3GoTiMRllFDGn1BaeWNfO6S0p7Cu4y4Fxe4kfy6dyU/Sm1aQ1
TpyOILpEKFxXRQHLWaIUVHvMGsoXmJW7Umh7y0Ws+nzLSAlCUMn3myuzhhGayXQL3GFInHHoo+Pr
SjsqcKhc29094ohXBt6u+qSNphwM6gas+3+frdIKhhP5Sk/ahVwQkuPSocMI2cD8JkS7CeDe4gwo
MqmVe2z/h5Qn7Uaz7w43hA6naOBg1+6BINAqnpSxODg6aRnAAJpPxf0CIjqR33x0blckwRMtAwMm
1gNrNl6PFlhygWlKYo2lmxGRV1BI9TkcdLssa6yQQSbYDUDyePDiNZOhgbm9FujnrNiERPn1Mp0O
+8vUBMwUKAd/9yGDh/JcaMm3xEL5ZejpmLQCyZ7LYdtT5jeKqYUt6sXP4MtD+s5fNtOkWX34kjuo
QxVQc8e64IjKL1MF3ApJb0t/S2BMI1vUjTJTCTutbSvJcxJ/gcBPPhZsXHf9RTskDj8a3q/7wpVm
CpwLjIvLOWW3sv+7Kb0qR4PgozYkF0ABgUEDgJcVhWU/SXXcDF/yrNTXpAZdyQ3x9BuRUf112tsE
AFB0+pNWr7stpPYMwYi+sl8rvPithMkiEd0vubQ5/2IP084X08KYChVjoMUATuLR56fCiXZCmy9O
1c7DNGj3qQXmLfywaQ5xrUqfPj1I/q7mcZWcQk2MWj2rZqIY+KzUXXveTxeRVOvG3OjCcXznf1Xf
HyOMdjWtgLzayjEqW/VBfJTeN8zyGRN0eA9nObktddsA5gKq58CN/fCRwOEY3pvoGmKi4b/EX4IL
NjUMC384YhUKIek2wayeqo9wLkhFwsIB2ifApDf9NZQMElfXBdRov9jHk5SQhKQiz3rEAqi7m09w
bKAcGQZLDcqqdwiw29K1kjODw+/HUlf/+SUwjsmzhZBOb6SDWr4PrpY1p3nL2Ct7tGcXT2e5lv7r
mnGH79Fh7ly3jWvziy8I9nIEHRsvpA9/BCrFlFxqxH1Njx8iLduhvbD6VIqgyLeqATWQ2i5XSmVB
+bSq8raTHoLSjkGiiZqMeHxo9GTQmni9r+uoJ4R+KuI7F/e0W3jsTGR65qw7Q0epYlZ9/SpUntze
ZaKXIz2DE+rsQyo117tpTaSyDbDWvDTwGEK4tReKHqecoQVOTyl8I+Y3bSfulLm6V2BuYt/hXB5x
sO88mrknxkHxgbTdpOt/ExwR9SQx0S6qxFenpSRMIIgE3sVmLewfzTjhwnqn6My6NHssFKA/1WLn
xkBONnLONCC1FpezNU1LimQBZP4O9BYj5fLB+i6K4HeCFgmerTDi/FrCM6fXYdLUi9vatzydHAR4
FNX/27corQzhlsgOn0DXktiRtLB1VTx12AaNItPXR4IStPwQ+nlO2XeJ6eLwZI7MXjX4lK/JxO28
jNfIzxFpBXYTQvBhJnbFxiv5XlAV+nephRL35WKmCyYA5CK7F4LhCurXsjXPUHJWgps2Jf0217xY
Uo6YB2HXm2q6lEZGwJONn9yfeuzl+vEeFbxN/ftyMQPxQJSDnrAmnsYU0sk8Nxg5rASnvrtLC5X8
zz/mdup14vIZvVs9Pj+ezhVSPUF8nFgBglhfC8ZOBY4P86KY1P3c5FOK86RukCxZEIp3dC3aEh0i
OFUuCtpc3XERIZd4Y/1R73ItlvQgYL255oi9iQSLdBjLn812KRpZbrHcAzpHrwFS5mmuTaiBmQs1
6vbbPoYz9FrDWnvp3fX1c4mB7UfGh1eQ0FbHqbAccWSqxCfvESyyjgfhVSICslFPe+98ENjl04Wu
am9GbGRw75g3n/k+ASADOh3mynABW8l5K1PAeLkXqcvo0BDiHMR9D5Rc/1z4Jc6qmsHwvrvQuDbh
1sP3+3n+C8xp+q30BIrl/3ynuPd+f5hoor0l4Q58wjI0xFLI5aeOMGOgARVcDwa65bZUY1r7rRqG
bV/zJRPfbi/jafof8P7tlhjDne/9R/8LQrY4I/rmQEJPpOieDmRbd1pk3ul1kYlgXHaz977P/K+x
xNaFKADNQesfS6GuQXekYGYmPErtL+9Oo9aqzewfKXOZ32w2JM2z905TMw3HmCuLhxYBOa8kjNBD
UASl6qZMBXnunaYaV7RZoxLtznUDGhpmj1+tpB6CskORvb7NQqXEdhjkAVgnFAW6D3LefEfgMaXv
TsUGa7yjx/RCI7pdB84tJ2nnIZSpKwC8kd6DrgS45i+jZ4AFKmbzb+wKw/y0uMLDTl5MM6qMwkD3
osTYFUIOKlPdSvFY6cttPXx12DHxIfQ2nS4CvPB2jqksiaoJ25gqQmtl44hXX1WoatXFxYRhRaro
ZwijZJBAsYIYNsmpNoebUXb7YAt9bG5qn/59ym4PIeTaEyz4gX6Sc5t+CTiYjWLLKhu/M8Zi5lG9
AU8Jfq46/NkVpQCgw77VmlKwijHqLWXKTbgANkt2zZ75dOMgDUwAOXBx7Z2/yNPG9mnSQCr5Ebjq
1FCF/cElEhjDsfxuhiwgIRoVKaA5iyrVztH5ang7T5QTmbN2BM636AFMFuOKjPBjERURKdIEh1pv
vAq8Bx3CD5n4LlOrnZnaEEKjgPb4ZS5hQAuVb6+2ZHGx0UyxYp6Vvp53bh+Wp3TWDRaZlbJkZ1X5
lJyIcRSCDuRuF+V7LeFvj0kge82XmeqoeHss7LqglpgY0WYmgDtgB5wd3M3j6MPIrMNxe72L97r1
s3DO7Xa8Y4wptVmzLUH2ZS0aMCVZ3BGLvJ6IDNu3Q7GDiVCkqC/6rAGE2/mtp0wWT7v1/rUD8MJk
pPDh3mykCOAR43VBCKa7CXkS6ONF6Xlh2m5hLiCUZFR1z/PLMrdR9IGEKneiJGDjuK7TnLP8R4hv
QOTRMu/EeXhDswlJ1LhesURIcBWsaFtaPEIeMRQLHwUUpnREpa/mE25HBv90AbIBfYL5yNS37Ttn
icLcGxjGY01IcOsv+ALVvz85BB4a12RPT5NiSNAkytA3x1PReMYKx5xx+PxK3C/myzlXByc+6+kI
a9RGq0Ja4pcQLiQ1pzLkKxnF48Yjc3ePMLWP0tsllnCBEd4TZoowQo0hqBv7/8gl4OmmuoZUmzAf
BrgFxoYaHmyI0CA/Qkzf/vAqZ3iD77tk4hw24wYFpq6/kYjZ8mV7niDqmt+kSLHJ8CwDbnOTPGmx
fy+RPeXHjCEhhvLQr1e6iTinB1nzxv2o39NE08ntWhhKag9UwvDKfomk7dzs9n8aG8UT3NbC6Oo9
UHibpYiCty1Wkz9wJtJ4jYvSBuy68dnLXjn8BLP2k1H2XNr2y2cbp2vUaujMUE+J/654+DG0aDkE
QPI4Rc+Ob7938p4Ow/OagdTDztBkfZSD9JyCCgoXU6eUcncd6Mc8ReGd0pjRDRS1DG2Nqd4Srzfr
Mwi0gjA/s1PEielCU/5XmOILjQKgD9/fGAvNSeqgXJhQauWhZvPAt+tHOUNUnXrrSd5ZKU/PToLG
SmzJ2YMSRHtmig4AzDYkxYtRfBDphI+WMsse3SYNC7Th1AVylJThuLBbZhCASPvSiqiTOfZFEOWN
T/F2dYWERPA52IVOfwnNITj1ovGv5YFE7troybvwIPMS8haUBGMJI0N81Gh4uRDnt+cjomzbDIBI
oJjLnP67YsIGKi8/euhUTr+8Ufx3LngSAzkIKiFLE++R87HcOgxheRKj/LWMGIyOHFh5rZpoO4/u
+POrr8dmaZE2HZ5yoPSQAi8QGbXNqGSi5LcvXHGEwyaXz7v8PxHnttU4GopPE3qsVZoxRoNnM+aj
jllVaspCYww9o/lmckhQ3sugD7JYs/hk8uJK+WK4vmDyFtbzbv2C5bbbgIu3asY8eS4VT4O5IZVg
JLA8/R7slg058c+eKKeay+YBn8b6zDRqAc/9DpFj2yYaAjVcDwUxY+18ksyPH7Lugn6r2Z/lVlTQ
Ed61RkoHBJpVEsQbwuc7yVg0pBVnLCt+sQbYw7KNB0zKz2qFyZtA/9rBu4qziZ9Hv65OcMV5Grsn
DkgHGsTuwb1tY0fktNNkeOh1rDFRsnADnhfIvqzk/r4CKYryReAWmz1o4pM++7FooUOagb5YtXli
xs4WlxbnpWA/OcS89kJrx1hIqgW/G4wqQ+rufiKqSMGGama80f/9ylNOfcgspBDpR/LbMoeHN1M2
0Snk2dT1Pe26TRhsm7IYKxb6UfOVL1Fgv80WSv7MfEsYRuFodZo8pncM9RGxZgHqjeixOrBUh/Le
bmW9aBDaAqJ3HENa9Ha+uv5jPtE9O+S1RmK/mCt8gIoFm3U9UORl6AWNqWGOlmr+GuEavyn4rDio
t7rEIpBnYMPy8gQjJyhSaUxBe9NtAXAHHWrznAWuv9+RXvrthkrRkGxkxUpckGhiitjmf3ieQs2y
FfeZ31rm8zJCTHWZVGmBV1rCa7t7DE/aZPh7nd2OwaTAoHF6SwLFjZmAN93GtY8OvWfPfUc4eo7+
6ZkgxbKMdbIzWoMkTThFvE47ggLH6so8nIlF3LxCA9zeRGkQ9wMb9rw1Nv+nxMNId4IhGpIhQmnf
ULmXP2ug2SweLpwEy0QEUDwKTWf6HYt5/SWPyxXwF7p1+mS7t+3PTDx7iDSP5Oc0E6Dra2X68Klm
W9Sr4kWyRJnIxQv6QkaLATyQlLZ/rcH9XuoZs5JG3oTcoZCDHZc6tEXYyhQWRExin/8jjIY9TZzp
GQEtv69aliTZDVLwarqajTZoTiLP7B1N9b20eYYEeZbxmzr1VItBJMksM0lIT45k5+L1zwlomF8b
lp7nadDVOnwnT0h/JN98kpYHIzAhRkhrURc2TO90J251y04P2wyPMQ56IoCOyzmsCTtZaY4XZ8Ob
fty7amxYx+KoOHlKvwf66hZOUu+Ojo5lVh4BKvZoMur06HWokZb4O805V9/wHxd/BdNNGJsmqWWQ
A/UJVKrOetVYfS+ODA0Chwu3iKi1hLLCSniQt3zHNw9lvUyNLKWp1YYBmce4Me3348uLpKNrlZ/P
IYLI4gnohp9kTiu9GNLfq2e/xrxnWwegDa3SjNLwmY56GRX3ysNyIGLC8XSpKBeU9Y7R/0pVsdr/
CseLBe3lw+MqClNotYmuNelNxLJHUA8vnv6rCAYUajVTGZMffXBwpaPatCAsxjMomjNxeQWWR4bK
aYM37wYfFFLIMxF54MBw2gy0xKQjOGv1z70Hnmxx/GNRafH4Ep/wjqJZYnzlG9c9zg/qObdV1Bql
TCfJHHyAb4/BBF/UsKiJkQKAPqKdBM3Yqj34kfXbtGfo0NBzd3Bv4gFWZAPRhqUSgUSvx5GyctIF
KEZd6lMM3xNE9BnuHiV0ebnDXQTJlslyIeMmaig3VRYccRcFBQTwi8STPndPqvfmEHo2LmqVMMzs
864xPD/q+LNuCh0WXSQgFgGfRvXzwRpgrjGnQ/XtJqaUtV1HzuqTsrEOcrQbbyze8Nbv618W/yo6
2LDdorvhvAnsepGlLmMVJ6BejnA0jpzIGPzfJCOtTr5WMYUz7eNBUICBkxivve2HOnxx0UhP3/SS
qhNfYtlC350zo4u210javbczsiFhBkdbSN1P2tnfPnR3gRu/ZGanX9ax85dHl2cB+zBwI3Hvq75w
FMKc0FaX6zorSty3iY0x5Y2bYDCAuIc6BnBWzCl0D+x2eMCJcf1CxcWhRJEX63sDTQ/O8F5ZvG36
1CyUhhzMHkbC5NuvvVT4Q6GSJQerQL+ltJIaKxuQYSnNEAKAa6COFt7oa8VffDS2Uf3BPwib197j
+u7FB0/jyC1LS9+3o89TNHGBZoaThIgh8bDnoNh3Zor2L10OgQ2tcVF67oK5TUnC9wjq8TS9P84j
xrhkNMQxLA7SbFgnc9NHY4sEYZ59Vn1xaFB5+DM6JrQlTajG2y8QoKJVrbyDR2DdKSeiUXZvHM7F
jrvi7jVozNictfpV1MOBn/wxvEN/kaXlQD8bL46tlE1VOFmaOQOEY8NRVEcs6W1W6uWLxBEZsd0V
uSqS12cDCIg8XK9S59GZ4it45KX/QB5XxpF9xT+2QhcZHzKfi+AvQdkgdk/1Y0BraLTH/dXrKj5V
u1oloexX44N49AlCmwtGDywVJwQxi/WVePg2DBbEGdf2mGUi+D0aF/au+ziEQtBvfu3SSevP1Waj
aE5eqkveX/p/Gt1ejMq0sRXVMSD9FVFSxoOzOhp/u87HCuXvHWTvzzhRH+aB2dJXkzQE1vChJQif
/zNTBxfQ6ndemWS77aWMaTBy7dua/Ow2rSsJl42GHWAP+kN5Qx7UGI6u8LxBMMwaCEs7GTH+QfyC
ap5j3oMFqJHLDwjWmUA0PLdU1cJckpQaNu2FkuYNlsUXPUwNBGoqwN13e066fA1UGzwSxo9nQexs
zUDuY0+CBIyRzI3okz2tKpOV0B6Ig56Ax5XAyyzJIEyf38WFLP+OnkmGzNWNiMVqnknsjtTZTVpp
YgtCSdGhDq90wZ7MnSmExv8jttfJANWom1kWShosatayaf2l9t1EafjwTGJ0TuElpGycaLT1beyg
nnMSjXF51zWPbdL9zHtKINaQt/X2nGUd09kdxX7ZUhHTKU2q4zFi7L1eH7wd4ffMWUo8igIx9C74
sqbBYgtn8D4HV9z7ZZW+ZuMaVmD/I1yooyF6bl7jj4OKAoWn3ZjEEjmFLG/hpi727sR/J6KMLZEB
xAATQORRXDBcUdlRkLyQpzzWkWkTHIIzBih1NbeeaN1Hk2nRr2mK27BELK329uPaxm76sBiD/HhS
jMHQuLxTVcB1CPAjozIHwhtab8kjzlEFHVtFno3w/XLYexL2Z9l+FyMtwdIzAM03JN6jssLh14pF
+uaCIJcAG5ct+SLbgL7QILMvBOEIrvb78cx5YvFqpgYU9gbrg5ZDDHlpQE8LVbGeMMjy7wL9sz3z
6QIqeIksUW/vq/8Pr+u3cLtGTCtYPHrThXp2j5ryo0hvlFIfDLQstFnTpOdc4fCVfC7F4Udf7f15
eGDogA3fV8OoEzmRT+6/bCh47xHL9n9622pSPyDaIg1TIj7ASj2lSr4J2RVXsqNTLDTHu7JtRmHj
F/uisVGimSv9c8heoA4icGml5p1FcA4Vdh67yAnqnEFrXKXJHK5Bw7EyGZlDgUTXkXNMdAwmd3gy
SWm5tBKrkoYt9Y00KgsgkR4gnSS//sbAACHpVUGKfU+iJwMbeCvcqRJvsZw/yBH9o9MEs0PFLs5W
ZYk/occdMZsApcjwLeCLXpYnfJD+2iPCC6LcO/ee6O07uCa6v41RYkGSV5w+cK8Fv6TTd4mpIrDF
cqZ7LJdMCaoJNvctq8IfSgocg98HLEdBo23Pcz5LbFcYtRfF0cTO8SnETpgb6yTMbUZTRF++R+1l
zwfeek6s2WIGQEYpiiEldPDAwAzu10kgApv3rVj2J1Eta/hxNv82i0ycjr1lWkYKFuTrxrTwrHgQ
gQOONKsDv523PV6s+pqHdIX0fase4TCatUMelZ+1z2tTxWUkDGlNeC958Rr3+2IcXnpcpBNywm9x
GbHeb0/6fpT/l/HXe3ZBofdxUYE1pl/m83AP6TdIUnXN5vd0aYC+uVYaFOGYVfoYUwXo2T0nAR+o
ejq3qRReKGbqQlTX3FDygKsLywxQ7AD0di/t/TSU7cFJIddpSmXTdR1uRRd57UP/FyAKxnmDcbjF
1SlrMQLkIEQ6FLE8KIivLzOMPVOjp9YovmPPHE6Gt0SScU5CMMB4ce2XH0XXQ6Hu8edf7wihxEue
TceNJPx55OeheZLvFpqZBOAO227TXpmFAcZsaRBGZZ1qy9hzG9WW+EcD9rpOjYRpeHUfdwysGLcT
V3+N2GA8NUTJ5S4MD3K75+xBySFH5yraCPRsLxQVjf0IQGX3W8rUYiwERA85mCrYgIXLWCJPXNYi
wLVCqoHpJsYfee2HEIYTMXSp63JhUFzgOeCG89qujVkS7EPbPila4l0KTVqYVBxA31OKol1mK/+M
eXPoPhkrlBwgj/srKuTADirsXgZbUOryQTQMzqKHEJNQPb8saLw6CwUb9E7Frxran12ZgUefwDOL
4n4T0pX91xNpn7OIKJLN1DUxf63lJYw/OnGEvSQKChvU4GfBsrmohRes0Ojc7/D2cGVLrWuupgiN
ziS1hVcxZhgFNR2MdD0HmlIhouQwq2l+qtTnF9nfDcu0wc5tMa1os8XYq6WVKV14csizzIr0ngF8
vAYctkC6z3111SdtRtTvWsuE2z/2+HlqZSenE4l5N1vi94liV0DLtSD7jeta3BsdEigmxQLipNMD
30jKUC4KGK9EupUmMYuFWZNthgUgLlNnFeQjuDE2atEogMuO7d2Dw7b9iq9h4NTPKK/9oXup2i3I
/88tiIBzB3lNOXyIBcoimCt0bpo40f12o1L1y6im0Vkled30HXXsS/I2aU2ExTCTEFnPLRDwc931
LlhNuuoPxCBP7n5monat7+vbOZHKf1ToxbPzBdf282mWqKNMQsvsVsjkVlrr8ehGrJvTHHiiT+jh
bdrqSurcgk3Kv9NnMjq7OYLIWI+7QQqzMOTbStZhALkRUjA+3EGYjt3dwgdsl3waDjuS67/i9SnK
xmMHqkLR8nTycZEhuvbq/ISkVj56VDK5YL/uaF4weKqmqz7U42j9dg0eKOT6isWnCx9fu/iupemv
REIfkZrNGahUY2c56hXCyLDDfM4IN/KPfUOdPXj6iyux7fVVNy7nbGi8QIpBXdu8ZqJatIgRr4LD
J4eL/DA3IUG/sxUmHFEvPOs5aMJC2xjfeGqf1X7ombPAAiJpc0mwVtlywENDgTTweaxCZ+7p44oI
3vQd4mv833Z57IyblBDEMiN7OLRoM0lAH+ptDBZyx8ghEE2bpJgYHSWgxWIeN8OZIku1Ku8CFInb
M2jmmj+jSv++6I5/SGssLrxQ9Hq7RMhf+lsDpyDq+pGMqz+Hdg6ArRldRaM5FRF/XOax2tQNi+DL
rPnpWFEqqtPP1mSOs+vwRdHfqCQrw3xOWPxNSfdzluluBwQU5p/V1OexlyPNckGteoBScPkMLLaD
LG27QuF2rKvRZTxpAD0+IUOFLPxZuwZs+dDc9bKA6IQjnBNdJ2xAM56c4JMmcb7IYH9YpR61QwyQ
g7M6ORAYFxxC2a1aUnErwOGxkiFP9tzUNPwBlaAwANtrENeofVZUiMm1k82IjyLwFaeK3IOXiJTL
dAUedvqwWRtVmztQSDrp2mXloxDfmdRJspVomicERqrDVg4ZRbmpuEP9kl12MnrlyU1lCg/afjCe
uogTlHNxGEko1JxZYgj2shQMyqloWBbRZJAtZtRcU0Ky/L9p/vvp/agBpib1b7RyQKcCYJmDkJmr
Lybo8fzi1BT1FQjncfV0JMucvPA+EHWBbUHM/hjIO5fw6lK58EMHm/jS0o+NV3VPHvvX+1zIh1sI
DlDWXtK5feDbzKUe4VekHs9bNYwxKB2r7qrX3WOiQL6u6yOz/amZljGocoH1heWCS9XmJkIHmmbI
7AGjUPtZYmQVuJpBYNOs4wfGCFYEWqLSrNSZSmgINoOiKQp1Dm37vp2FB8Uv3LYg6HvnzuYSrQlN
X8yr7tLB5He8hb/GSHcrcH04g0ps8/v/U6BA4hBTSuKu3PUMG6VgmChtwzWp9tB+nyO7bcTg+KWs
CazkA0+vUNkuI6qW3+RvHX31r0RkVnqydJDHdewMPfBtVEvtVIeED0JqrO2r9hAQ4DUY0xpJaNPF
f3tyXilttd0dm51Uyrn/4iYirWWUWhy82AenppI4rgWY7/QFcczG+ennMFpremwgc9RoRm3eDJTi
kTJ/1Dw+GzN6/03JJPP5oBFGuki8fmKzKHaofM/sC5inNAda2+9yjBVuScg2QR9npPOSnWMUg06g
wGNxFzzRwdxA6DPY0xHi1AqrZdfIMUI9DW58pfJm6Off1dD7oc07RiLvRouWo0ucKGoGmW1kh2Mj
Ou/5WjI7UIFwHBGJQ6B9dqQJpPdeEK6RcgSw9KlbHjwyV/E/nUti05ocnyJUpm7xIp+b++uXsgEF
d0cjA9lhKHrdfi7p4rFVLqzJkDoidSw2HvbIwzi2ZPwwdN+kIh0k+XlYN4FrBXLLxFokvIrVkveX
iaf04m1YzBBJ8q7UdAFJpfG35EkvJPHXkKyimNhIgzuT6+Hdn20hffhljx/6MZ4MP/aXXu2DgBXc
6JP1q2w4EZOw/PjK1LtnioRPdw9RuUmGHMrH+Xx1UvuAl/F0guVhUho+cFicCxJWkg6O20ssejSd
PmMxpfSSDivzYvmbdQ79GtDVfM+ZCrTRobt4lD9+tU4tSz+EfxJhHKdXrhpV0Trs4jfCCGOQsX1k
+kaIfr4NdMtxioHKSLmZSTXjiwbODGkEjtkaHBa7VHD4FEhXOzLuL403dAvUVHeSYhvbReeJWeAe
EjOf3Dk+mgxcVpKO+ZsAhrcK7vEG85V9/xC+IJOzmZ7TyRHOmzTp4Ky1+TAQSYorjPBryO4JnGlm
vzD7fJuLI3r0vm041OBumETIs+K9x4PYBLzmZ7Y7g5Msx098YUXWa/R627hdIPWu/6C18PRsMD16
YNxtaPQHmzbIjQAzGSgc3nlewumFv9k9lS9wgcXbRg28uGGXaANDAcWRk18JBLAYO6oP2lLMJ4Y0
uXYYKgji/IOXMRCwXtAtoiuqRFrp2AINbd3PE/SZ1IwrMK+53cviREZic797xuHNokY7fXk5nRlo
eDQBjZMnfe8bvBcc4FboxUSJeI82Xb+PejwMOOBwwHD3mDa6cRuYHGpu72X/fjoemceyoi05xzgQ
145BoakDPU2KL1Qmasl29BYZEzE2QytbEtbjrQipxiPP4039Y3H2Y9mPF/tPoIzxysZlJUsQ7Zpx
xygnFMLfGQUMxelRfrPYGRlLZtG8E2+uQDS0xk5UqBh89SYlqkVqzseUdSQJnZc8YOei+BogLP7C
9vdISppL+sX1YagPmPVvdw0lAJRPgglbdVyrbD1Qiqo9O6tdZfDpNNBl7tRtSi7cteqaIjK1Zmt3
pt04Oul6G32EjQyQiISq9pi9bZ4oNOO4RPnQ9U6+wdFtAzVE8MPbiImWJgq2vS5lCl6b6a95JZgp
Glc+WO96kLXxkQGpF5MTYFKsYJGKzelPOYsCSOUSk4T463lsclZwXeirNIkvyPegL0g+e4WXuUsp
FJQYeh3c/gBz3XFbTuNLSrvzas8lvIVHaLgwwdJMdIMqBSbw/RckodJiNjdb/TcM5jk6/Max6Syf
Pw4i3Zfdm6PbEd7T2fkRaVu+tuLEqF79zr/YpsreGkhjHnC5GifpPTPMVjiF2ZvZpViBvZhz3o1p
Vj38URy6xGrSKkQujqH0N9xTKs4gi7yG0N2szfKTYlPMI6+Lau5KzUwsKj+V8SyoozgjzeoZy5ue
wA7hjTirTSkn8vYUkgFp/aX3dg06M7W92Qs5xBmKJs6GNGkfLbu7bG5PZ8pst7KjR/m/n4vQS0BL
/VUhmz8UF+O77P8TOMfIGc6qN4C0P9BYJoAiSHXmKi74pOcX0dwGKJ9PN/XOSut8e9LIrqmX9SiH
OCVbYdu9zZSaIJZzoOOVJzj58Ik618/nqvuoE62z+/yHwj1XS8o2bhluOQj49I6GA7ILk5nxlUpg
c+YW00/ozSWl9slUNkXpVa2KmFLslPBgQO0bHBXpv7/fjJK5KA9J6MHihi24uyb/8wOdiFElFJL2
dPEYDjMozB+UCWLtvGvfhGNfxQOURduLlqbzOwWKRCZGoQ+Cqo5oHoxaurJ4HvsfeoSTpExhz64q
yo1J/YT/fF6TqTzrtp2tlZGxMsedbGQ8NtgZNg6DE21C2zWbmzlcUUwUn9gV8pllOrsrt5UF3RVN
o0PTeHV7AKeyFLm5zvlqA2QijZ+2dFFtp6AipaaSYl6/fb+uBAQYS5e3ncQmpL13eSX1Hn48d6To
MNOeZIpbwKJSzONpaseBC3ZVd/5q4Gc32hRVs+j36dmeas2+WaIe/rfd/j/y1ySGn/vzinBOnvYm
jBvObZePr1cd0aqZFw4cC/qCpNDfShDJoUFlmBzDdLc8CFI2CcgfJAGllZwt6NalOFjZdypSKXKQ
qX54j/po9fkfXV/5E8XgpDHSDhkENRu+lXlMlxxLKg9xL5O7Cyma4TLb9R1O8R1nyIly7EbD+6CL
Fn1BYo3Aph9JMiulOy5k/fj2OZU+BzX++884YiITWyStd2JaglKnmSapCn4zNAVw3QB9qmu5SRn2
IQJtVZc3AHTP0dJjL7VOMuKbDq0zIWfW3U2SE9NGtvoBNEDct5K21O3pVqPCMxUz+XicajnUKwhy
So8MghFRtcvLKLc5ksSDQgUlLtHmWbAwq4lEPyMf1j2u/4Z+Uwj4EBVr0U1x5rIqq9Qwf3NOKXOt
jnu5T2UG2pS1b1LTTpYikDlTb/6iW7ZHu+aNqREIb7eAWt7MjzKWVUPEbKsLvTceSYNyUQKVqGmI
DDn9/Pc6k4kI3uJj4clX9rZjfpDRllkmbSWdiAFmGu3S8QrimQxcMa+iDovpBiNso8SMmH61FlZU
llONUbPhu51oeuBnuPgQTeOG2wMdVrmOM1ftSELP3sySwEZAmrQ8nDCltNU4aHooIfq94ysfPfWA
5gFyB7ybsr8+3eMVv5HJ7CJ3zYE5iClZO9yCvE/G/uYsFVo4S2HjxI9Befbz5igU05knwMFljonq
cL+8ylkV54e6m42TLE8X5qniGrlDVQpgEYVdNmgnSQmnq3aW8Gk1M0L+p7Pk741QZke2thbRUMS6
Y9TeicLkV/hDwnQ+epfOROBN9zIZ/dIFCXHVS/cYpgqoBPhjUf85CGEi2Ooxzp2PY2E4uRYikRIa
TfUCkyM4nQ74ZWvcMg0N02qxf3hNVbzxUtJiky+cYjgenN8UYAm1xpSMvFCvvoDy2SaRqK8FJcSy
c1s+OX97ubKTBBEuNLAC88jnhYf+CN0LFKP5aHB8nxTx+8wz5K6w9jWBZDQTkh+YDG/ILjfPL5SA
Ac5rbN6g6Aga90lVpmIbMiQ1uBRPBHGkuPL59FzL6C105qUMj1HrceSomQFm5LGvgBYvdc49ypeU
ZvoXJ1HsQJVm3Uzu0LLUlHdxlGOoaq1pVYxN1IZ35DQgYejIximFqDbKT4F9HQoW6rwcYyAUKcX7
UFB9BMdzrWQN3BSjjQ8dq0wdat8Xy0siFxLVgu204hzfFySgi6vuX0tlKSbKrqY1nlPAr7Wb+ZLF
RIaI1YT/cRMTg5HeqtqKAypgHPVDuL9nbBs4w5owrKKev9BDOYEEMDs9u1F9lAQn6Gmyxu3qbkA8
s47mCPHNrEG1wDrPDtaLUVhpdwVm0I01PMynLf6xzDHeCYGYp5ob9Ez967Cq8DVjHM0KN4GY5Twl
lZH1tM26KlD79S+jFBJ8iQGnftpudkf/AVXvtXJBknrfiKpTKOwmK5ma36zYL408iCA1i8b4ODbZ
ON9370AfCx41De9Trr2OmTO6Oo5ROEBFx4tvuYeHxQtLm+aKVl8hzQ19IXV4jVbzrcRjN8uDk/Se
FV1QShhTuUCd6pcvM6hfaqdXmKtU9MfLQV2BrcDXv+v/zAhh161/r3R9hfW9VLD4vRDH8IiahScl
OvScCD2TOtapN5gjrAEN7XWulQ1jh+GL5BYITisLtURXpFu+6FYpCQhwZt143XgH9JcHvvX9zOul
moJmfcZd/ZzBfbGy6NtOoxLyGoLQk5up1yTSjNk9+niWJCEeLepxo0LsA+Ye9EAOqp475Oilrpp4
w17r1Zig7HbyBDjGZZHIHCdO/veD9ZEenvnDQ4cR15lBCYpUBGS4Y8Tysp8dywPLHaG+RrrF60cG
ZSGDpmfhmYvBJMj8SELnnk9PUfz3PRU8Eq9bKWFOIdjqiP87I/Y7GjHavI8JyWvP0n4SGrBuZdCI
ACzwdc8H9qMIwaIoRv5P+JRQUdSYJiiq4faYleYXo34BliLGWAGFk51r1oGsbtxWVMbxhcH45+ZV
sXN1raZxhLPyV6OXqpkjZuU0No6ZPvWTdd8itSdhXOUkXossYsmy2cdZhlIyxC7+Gbi1GouEDkbJ
DukVojL/sZhLJvMfRS5qpzlmnzjIBgdTkM9+YGa83g7Ifk5yq/jQqlLjR8JG2TgDKAKeWV4khf2b
o6UuWLCb6pq1sGYeAvdWfYzp96A239EW6nYh6DXMR+yfeROrtXSc+uhG2YHurlWckVqIdHhgKAL7
cDHA5cMNG/dshP8OBHl7w4sx5lxkHLfaXglzxpJELO4YA/r5fOh1gqhj8FbEY2aGpSsQv4PRm7Bo
G5D3Z8MOaKtFukVvM8JjZC3M/76DYkO30WAN5yOUFnwOhMMKYxCLaJI5L5+jXWd38tLUodZv3rZ/
Gx/h4fflfAX/S/1z3jIk4x6hUMx4U5HiOnE4sUbVsKPbNbojdXxPkIy6vtWreAHqGcOZM1+QZXZf
YuihYlG7Rf74jV1uRo/7jFB5MIaivgo8hLmyIUDQbLkXGpJHZb6IhEPLTpFJVUCwv3/nB0zcYbq0
IZnWGFluHBDOkxdEw1ieI8+zF9zlDR4KC2k0z/G9Dn5979yCICSnMwJXXA6bHGVcrjyuDdJgYfRH
ifHEmI8DxF58YeKrhjLG5NevMAgrocZtySxOjpeGhL5BKk1PpSWQTCsHw/RMjhkZUxtun70fZL18
a+xY9iYAV1DiJrPjto5aUdposNvDYy7IecEsfTK3gvTmSbo/c9aJg/pBWbngSref5skQMdANHwG6
SIoNWvkwoG903zr1WAbPRPIPHr0g0SCV2gswJnmYXSVS2WBRT9T1psbrs8A7oD/QUu+WvRsehC7x
BHSP2PQB0kpA7MXv3l+L2Zessrote4O5f8Agomuj702G/XOOPeiGs99BsaytW+NlcqUTGRBw/2FK
K66Y3eCihEnOIqpwu124yQuFV//wzLY9wHX5PftrViPFEvoNOzfODruO5H/Dh2qP1mbVg5XUu+u3
+EsY9awsRr9TtSJHkczPIwhnZ8dILiHHrFSGCO3Sie8HxKxGsb34vUA3bb7EiI/8w64+fVnrBoUV
xVBpGJVPyqs0CagkmCi+wcrVw1Xpyhr9hSykPaAbYElccff9anfseZ8yyoH5MiJ7UXxJG1qH7QrS
WeQzE2fiaTX4JlfOjMxD6ouaXwYEXcG/+0XIMqzdfgDVV38DyPAoNYbGOLMAYJAUGTRaF42tPUnr
9pGr/VrvN2qZAdQQJ4MhZ9qqkxzyy0rxMd8iCnl7shr//88ejRy2IFjw9vqAaBZZ2KZi8MPcD8Lw
vbC9o5UVHegC88hAQeTN2dS6gYGZ2aJqYRxx6Zjy1EZfXJLWDI842/Y3/BMTOQwRonh7lvKeReQ6
KZp8QEKxVTPZxlfrPq6dMRdNcwoRH2VQB9aHz2nLqi/6mzCQBm7b+AO9fJhdRDSavfyZ6ka2iD32
GIHZS9i+VYR6poUsBg+uhzTrtaHoHqGxfVtJ3FmlYToF/7wjGC4Up2QMgwdtnVEOLopeBfRAEgqK
EHJKB2GuA1I3BhyeeUJhiv7sdi7ZtDuheSuoI0KXk9lXdAqXyUoNtB3mwqoOQXOX1llchmhPIGAt
JhjdZhhsBgmPQ1feDw6c0pcjxcQDa7ceaIn3iJrhlyw9MAdB4+dKbHcTdlqNJgkLDBoWkanX77Er
zCiIexeAy455xLyBlqvTkQIYrG8zXljTSJyYmaiSP9GeM0gHXtLCdZ/4oJCktuWCb8uyPuuH278d
dm/Uiv7oc3DAD4xJdkV1ZwtCT4od4bawLx0sv4GVSSg7B6WnEPF5qYyQbnVmTCw8KjxFAiORuvEI
9F5s1VUEYNRcRlGEV+6758X2qExNb3GvHXUN3n6nq+eelorxZ99st3+5KnpMmGVKPJD0pTktaQ5m
rPnweyiCtjcjLX/KIlxFdBxMjgOwmnz5zj0YZxvH82SLrDYkah2xkLSKKg2akpITBRT68A8pfpD1
ECQ/WjQJM+JORDf9owUcG6KkFLpa+OLQUJnK7B1Pcz0KL/DMpk0p0TyCzRSmyZ+y6khGguny1PqM
323CxDzwN2ZikM+sm1tjZmuogfOCEnMyXiEzQl1wmbZCyauIQ/zrXHyiufOx8kmVAyMp1Slmj7SU
uHegJBfr62YerW9UmDf9PHu9TeSvDEV6P6p2Oh6OAE5U9eT1fD3VpZWpgGeSyBqwwxDKuycCXhAn
JcLbIZo52b6U/15CTh7/28YXen2Hv0Uo6TJ/OKMPdTQ4KKSpe25CAjQyvzl6VW8hI0CS6PBW9VxU
2QxxK34pfCm2uFcVPQWDFEwZeyJk2B+R9pcLrxuKlAkQ2KDsi0KeCGsKTIKrgXT4YMlyVdB1uGzN
eIeWXh/BRHY4nw/M4IzXJ+HOYufsPu0XZkkthXdeJwlf1P6gvDByHvzPz/3qytyzemGVsyhUYJeG
2FL+jeROzfNacfU2efUKJ+SO9NNY9WL1NN9KDuvd2P77SbdxWyJZayX7j/Qr7E1JMoi9IlYvAwuF
pxYwqOLblQ8oZVT17sPzMP0wJRguPWQwBq+skB8rJz6rcI0Tyl8eYx2Y08r6RCXUjEEu9RZ44cYS
REW9BeGtMkAeCz6MsIFcVeU0ehz9i+T9vP+dCUzh3pzIaFl3JM3WJsH9r/KytCT92hUZjO+GKblg
K0/6ErJ+Ea4ff5Mn1pNFQJ9pznYathwnWDnfEx+CSQXZpzL0AmlhNs3QKqGjg6q0FlaU//To5Bnt
MZrQGEecsIvniXkO+mQqdbOxWeF241b5HRUNXzlnIzYc3X5bc+x+miqep2/pf7aD0ziawnx4hjkJ
awIUN2kyP07hnEd1awzfWL3V4jz6OG6TzR8GeKiqG+1+LZ0aRZ6zVHuFwbLvnJjKruk9W+tooO4A
YyxV5uH8izZD/j2iDECeMKBhLvV7PlL7ozRT/QLHLmp89rbsugbu1zhGaJdIbYGGHsUqoU65sfkD
ot7cYPxn+soKnjWKPpubKUVBoeoI7WRzKfODy6C8GzbNixmAbmtCmncRbqarW1ReWlIbVQG0UssV
q5pEQkLtlv6x0CeA99iz/Xbk3PLVAuwjflno1aMb3Vc1TiAbR+8TZpvv6RJbtCxgN1gvpTF0bqPA
ddUU7w5f4vbSU3DLAp+5UxxQkhVouoNTorN8DfgBaJ2oYOO0jkxmnQBbSsGPS9em6vS8zRW9Ygaf
BqPeqKLLzB7JQKcVoR7CVnGuZD80WA5tycy5e7QJxyeG7m870H9N4hvK6HBB5MhFApVifGATRURw
ie3lH3rEVS6YV6rD0QR3eeZ8NikR5KzD6vqgCDcL1+/GMjXqHfIsGMkkak4ySpL+9tSRMJJ97SVD
fjjTVBWsTAe3BpBIs/4+xJUX7w8A58wzP3b/oI1jvzC/wB6IOlgsUHZXlJ32c+iJVNc4rAWaPfKg
JkQfJNpEhyxBgJ8JOIJZGRYemChtPSG95Y9unSlOeL2eml1nRRjNo87ikfdR0hw4wDq+Tw/Fdaaz
Xn4Qz51Oo59PbfXT54/PxIlLLzqzYfUUzxMrjCaKCTAi6ZX8DiN/K1G/Qqyy++tYiyVvxglhDEdM
geHZ33rJWOKhVnfd6O9hUxrIv6sNkWUyqcem8CEh7bpMNR1UdqoQZxBmbPV85s95CtT+IWAcgQIQ
3+ScYbjC5fiQOvfrqdohSdKi2Xu/benY2Zs/sSW/0aSocSqKBH03mX7h78/kiV22CC+MdBfbbmRT
M0Xh5pAq0MZSJN9+XqXd3i2NHgrqHZKFllpbtmnNBnLmolN7GXRK7T1wtAVdIJCYVz31Bp8JP3Tu
awdcvb39ARVvQYkYo5Xs11Qmm93DoJykTxpgLcFM6UDH1BYXrgK+4xT0ahYPIHkmk5h4z7QkAaqc
yNstXlpAAi8xN85XWVFM71NSpNJDexCxtURwy6JBM8KKzzpY6a0AiPzyqVKYaK0iGyE0/j+Spb+2
sD56khzq6jDJ35F+Mrb17FmkvMn4i5KhwpNKzKceKyHc2cfDfMXU/qDTvcbxbKe/Klpqb8WMI4d+
ovg/YtUxq6RzeiJD1KtMr+/kQhjrJ0KmGDPJePfPRhyYZLC4NZYDNIxDXKTijaMfRl3+SomSUFOv
d1Lnoy3PXFYAR4d9ZfoBU+9ROWhPN3BdGnBiJZ/ZTVEfp6MlGWxRQ33Ebqxr8P2OLAyO46VOK8zQ
n6SlsgAN5uWBk+OiqWA1bcTBxniaqUB1Ixbjrz0JUOwNZiEFLnLf9HVPhh+JnY+OBcu8iVSfhcAa
gmxYMJDQqL20cCn5Ep5kmFXWLefSKWKxPXILfNpbBXdpLoAZR49pew/TNKDx2vsaM0uXTnk7eJFq
eyStBPSOuY/XrUbMg56/xcLiDkJY0Wd1Ac4wWr1C9eYABmfq0fd/SaLIvl7b1SrDrMgW2X0kiAOy
zqnyZgC6vZpqXMdn9uCUlY9smegkqvCYJPAfD6l+43l4HiqKliWhJ0tnlGEmEVYCtfD/FQToZVak
KKmhYbxAUSVnMg62TJ7CxHhtA8aB2FBvsGhD1xGDyvnlNAyyRAebJxu3wxWIhScSF8FsK7YU9DA8
9n1xzMNmzIgq8ULPWdWIJq6xwlreoCY9vA9mPAbDORQEcNqRw+0AmynTI1ezFk4xIA/D63ALMIBV
julXy7tXN2fkShzwolgVSjssHjxNAgfVyoj92JFCv+IETPtiy8Yk2DU9pKVWWXYhxNxwPu9r0l/c
ABE9FmBa2eL5acOkeKxsZ13643ng3rHEXjtrCfMKLntWh+CGMvrDiLvaHfNgqAuQtw9FQNiinZdk
l/XkAYfp3qYObJq2xCVeFKaj02XR1YaYWlc2uTrQc7at5co7cqz0DYv3bPnjrJpeeyAKTOEud6gx
exrF1/3Mx8gCYTzEod+eoSqdHYxIrf+zp79I/B0QCGiuA1xjgo09FKlwMehYz+CqJxnYUIYoLWXo
CG8d5Hy2KLrg0aeQl5rzUS3waGvWXGpjvmMowiMuWMXuVgQHu5ozVkfW5moPb8OerF+FxdSwwtwG
wPiDXin5T5A0xB5PqXpr2xqwZGznhCbb+n7dQeHDdz9IE+czDZzoVB7tSq14UtUh3TujsyKfxddn
fYJpdsIm0q3ZnTqu4j824ZQ1mWAJtHI4Or6dbTDtNVRtojBu1rzIGPRm6CvQp+J81rWbfGH3FwPX
998H/fX3pMbrFcBKyxbQ2X/5qLxnmJHMn2cNpSLHgg55Gjocz39a2EEjcJOvCc7RMu4G5Z5Vf89t
NRLV2oAmG71xhYOcIp+RLOzwmS5eUW7xpeBUZcxs5O9B/ywAyupEAhfdqASDKzOw2SmlW6z9MXRy
rAZiYGXs4gp6dqHgrAKRNjRw3iq270pdq9BWHlR2SJjM2ba5X6YpIlOZ8i1Mwb9oL9E9PW0Be/Lf
Q99ejfnoz+1+tRx2c7lGeJBpaS8m18fnvraF49DcGadZNzaaX1fEV7CuE10BD9/SZc0DJkg61krb
OW1RxyZWh9N47tVdh7LG0tWLiOpRTJFhqKkVEBPwGxsK30Dbm+TWIOeIJUlQISf7+kUcJ22yXoPZ
9UHpsFzFW9l7nNS1HAxxStcm0NJ2bL5jVtiCsgFVdTo+Y/pjjbpF5ABS2VAKQV0lufueOpEA1tGf
hS2HyLaMo/SHxBEElC6UtHZbWXuIRi8owWmC9+afjFTayFr4RXpbB2w2lAHhyF0DppwZcqhV7R2O
3Zt/XzgbydyFvzNs9HT36UTwU1t4ENM1Yhtt6tXyL2ZAtayvK/QaQM0Bk53IOZdRUk0yI2f/I3Ry
pSJHtNr3PSFM5zrEgLQeLVidlGl/uURJPkN4mymWLuMeUo0cssb+EY7A5kNo5ZJZpFkfulo/BXAl
UC2dAnEj9WnxJ5I52QkRJX5xxBmiVW+HV358hDJFpnra0G5chEz2JIgDp01SjMptIDhLKF5Yx6QM
Udr5s3feGPkd2PvYePwk4oXnNV1nILdDMeupCRtex4jb9kGQnJuHoVvO7LRYtUupiN9lW0YK7iqg
ln6/6C1i5xSRX0Gmr++RCa5jsKqIFiAt3XikwRVlU6jNx23blm6Y//VisKM+SQ3ikqUSmaiHSj5G
0KfUuocGL7PcJrqNQ2Sqh7O7jeMahEXzgNULcJAZBXFrkzGV5ZyghMXzKF6nwI3p4/zv9yDOAoKP
jiSrgczGnxAX7drOMxO4xiMdLs/e8RuiFbxA+xrPmDJT87InZ1DP8p2ktyKOLEqpYajkm0wMgm/U
G+cv9I079xnk4MIKpIy7BwipT5teGH+XDAzdVss9Ul8dbhPpOTLJ6Xw/kcH0rl+7jBJhUFsLKZEq
6xCVHkbHTHl4KckErL+6V0l70NG9HdOvvkbFKFO3aBg8DEfFRlDqjbl2vBgvtfcYecQaKWRjTIbx
bXXwYxN/nNEGUYepKerrAqDuoJhrIvnOI3MuQxiI0uZR5QDM8pjzjaOQkA74MLtgXOOArPzFbDi0
RJhjMXCaMbgB7nZNItvBLntCixDDQTO6wJ1d11+o69JPtBtILkBC9rlnOWDkuuXktEG3h7Jri9L7
7jIEeHyRKydfay4vNtLyP6hFpc2xC2PuXpmxwPgNY0L1fe1veTZWxuSFIR+M38/wMTyCnLy+9O6K
vJFdmh8DQHfPpqP3ClOXMSQ9J/3zTG/dAzwTGNKfr6IAlUFK+Cl0lIP070bohQF5iyNexsyP4NUa
Jv61fH08KFXg5warghqc69ErJ/YphL+FcSf5xBFsxkF2l6/qj19z6geWLnqZM7D/HG9Kvuszbh+n
O7VcGogUep2vbSWXNQc3/DYSKwhkO8QTtC4BSRN0fVXxXo3T4KQlSVnKgmqfEG5nFRJiCgz4mlHC
FJGmIpAs908I9uYro4h5xzZO/vugXfRN2xfG4rkCeobSw3A1ARoAjR/cMkRMzH+HUvRbapvfzckh
jUYvAO9UuWJ1BCZcD5DW3k6tyGul24kACDCgnufHEOVSJ2e3KLbss7AWXJuZBFsivU2iQbgzSfIz
TH8/NHUZnQgJ/4oco5VBcotewJFq/6QbClb0ZHlkD8feYUicUUIar3lHoyRgoNF23sYQt/fssRTF
dz5yRy1OLqDsOzTo4rXbai7Mq0tQTRz2DEhMgvaVqGvzjGlNMN+JmWGaSMN9hEiEc3LhnmIyHEWN
C6XKAQAEjRfxYX8Dbkq5gqUZE4JGUYDr1DFQypJ9Tkpho6+ospzcZM/1Dc9OAdz8En0Sy9h5EGRO
LF4PQkS84UOQ6pnEhpYv6P39RtGSLuEqTjR3PpjNb0hwCjW8muYcUCzEr4kj+rMSjlf1V17GulJW
ij5aWQv7inLqySTZnXu7aLusEpS29SnT96j1oO/nttmMIvnGIiTRcQ1JUYaZvVovbhzKnErD3H8+
EPA//mjx9S3AfihSvP0U6Y9JE0ZFGlJ8HFioFNT3AeDDF7bP03VeDmyvoneV86IiBjipLZtz+409
c4qEX5nJ/sepxUyt9ocYDUMnlXMWRRnbnpjIQbY0vNXXxnvoK3/1tukldVO6YXWZdR5ywnSg46un
4JyNBMr2kMx/LLsiRv2QUP+GjYulaK4WChHle+g3oxezKMF1ftbHofthIAirGMJcUUWPzaSdKuv3
BhYJYgPhhO76Q6dWASZyXAwGA7Yf5PkN2qdVBpfYfGKitu0OWe/WwNilsKlNIAOiVeqK3nsqpx2v
k3/8j45O6Gt/Uy4Gx4UXkKUfREXYT0p1Kimdv1Ae277JlaUnOetC514lRlsyIYrInvdSneIb7DPv
j3w7foeld8sZZ+vyRjv4dltWf+omr9IhR94rJbHHAb0eGOJYsbj6a09WWAYqHAEAvp/03nd5iMc3
WhYEZCg/9zRtfYVCUq0SriwCpZDH23DuMNzpeMruKT1WT1BnLRDB9nXMdUzwwo2D7cUXKl67BuuH
ntPhB9YcKykBSfM2hXzK4VlOlFtlAMpnJvGFoRCDKydIsf9OzkxN6whXrAELMG96d41esrnUwQhl
1I29YBLp7zwqjQh4Q33qEuoP7FTrbDRYcm9FxSHdFw8jUYXq20e3DDYe56CR8x1OVjqTOk5FEPBG
dH/Oc/1cDvH+Nl8d/U1x3TFxWfxDp3GdZ5Dnxx/vhnxzA4BLiuCvphwytST76DS7EFiuQD8oA6a+
4cOD/y4BrI86SzTGICqQbTvoYp8hovOJ5QbbQLx6gJv0/xOTn4nXlX2nVNTlJNMQqoql5Ho5eXnN
bZZVyitlxNw8Qye0qFwqwer5bnQlMrQ7ewHpT38Jiskd5t96amoaYIf4wZ3HCCJZKAvPP2g7ZFyr
D3zQf/JzHEXP8h5Ym09Zeb4tLTqWe52h1ic1Dm0ZgvLMX98DaPDsZnB3Zx13hhcFWl+yA9fVXgNH
bIN2yFBhKbZ2zEQRGkbC32Y7aATEbAjKvcPb3c01diNQRzBWbLg8G4ASyP7z3T+6cZ1WDeRhM24p
FwuyA2KElKQh0AB5hVJt2DTDOwy8KJf5kztJSB/esTws0JzJ2uWBWqDqIsRs8pQDnYc91aCCDjUJ
dddTzc/QbvFIrtTuo5a6wINdEB3sLqceWnfhsTuu8bC9Y95aUSHzzblOyO8IGOoAFhagF6NBz9in
jx9Bcnv/dPQXZi03LnGoxybrXfvQTY7YggkhynSueeS6oPnSk3KeZFp9rI/Rsuxhjfhv/GIjG+Fi
jjAi9JaNEDylzmqCJKO+LUnq9z9ojFH7IYb1Y/tVQ7o5w9yJDkd636G99ibV4JmxQ+nc4Md1B0vS
rhfpW4x5JQ6chk37nqpA92RgkkMzOLp8/PPXuZP7HnGR01rr+LM2FTiShRtrhr6rnHJ8u8YHwkGP
5xePkXEDvGP5VTzXk6xZdNKhtZbl6bb4yNBd32ILh/R+nN2YNr1rKyENMzub54hF7qe8z51ppcgh
3B3ZNC61tFFKRDCPcq5W5NrucmJWT9tyN2YIGyTcAkdmsHGteN00izeJy73Bq8Qgo4K7kpjIuihb
vEjuKHW2T5DL+eF0R9yU1+Loc1Ctfl0JDzMYrRj7OrHAcMxQS2v7PR6kotNHo8xGfwXmE5w2ECKQ
xD7/3feCtTLr4L7lWwv9BGA57r/IL4UGgtVJ158RdxFFFZJkFf5Xiis1PN/OKlHKNSf+8w3ea6vP
cEsi432NYSYQ0myG2DEzHWI2DAhwmqWdmKh4pjbFFieZhZkG1Cf5nrREnoz7oTYCIfXEKiLNNvt8
KBW7y2fCkubvjElR4aPQ41jT7h3xtbv6kF0fr3AOttSeCV2qVL7rlHuH0g6axnxQw3Mbveyc3eG9
9d5kPENtdS0JO1gnpLYtYAay1mSy/68xVqMqURtXBA/Ushjlr8JVXSnukm0k1qW01iy8rbs8mN20
YrvSL5ziHKnby/wCcEJ+w3+5RMFLE3gZi0Lee/M4lKK8ryLZEfG9OqqGGt+kSeWLDmyzjvlyrY4o
2HI38OOseey2RiZ7W4tRLBqQgGYButJebBq2lnLSBsqVQpSibGKbyQeIkYAr9GEvCt2bnLWbBP9/
Eub5pDubji/yuH9DFG1hZN1+o+K5XNBSTSJ//hP6fAUfR+U7tFGjDVHi8xgaXuWq4187CJsvaKtk
QE0XTdSdT8XWCWjylCFL6+N7+tJJVWcjfYYl9uWioE3f+2sIZKlAZk1BPwNFflHlAsUQwbu9GhF5
ck+SUQeYnYILej8YGxqA1vFFkasFc50EInF8XQE8z61w7ZTtheu5czFy6B4+LTlpCard/yjn8sq4
xsS2p9YjEkhfU+0YBM9He2k817JGAvDFyFissTRB8V9BIZ345uBB09Anz1snDjcCjGL2/8m5Y89V
f4h9MWxx6RYP/MPrU2cYa+/VvKnqizuAAtrRiwj14V9K83tVNI3+pyEyqtwzNwmno3U9EvE2hTJg
S6CtLA4yDH8G+aKrEP51NEFxmR75XDdMn1S2OhdiQuysbAUgufIJPGeSWGfQEajL6Ru+cCU+CIpi
WIJL6978ZYzXppsjFFtoevQIRKvctukvJldBFDK2+K8GgFV2Ef0BRMTpF4zN+Ixe0kN48mKW+sii
TJW58lvKHwWiwezrZp0o9d8Q9dHTOd5K5fPG0pvXsUUnYEU27BOngZlClr+MJby3SMrAGdInEXOz
5HZya6CrXaRox4PBVCBCIaVo4EZcuUUlXXUEwje9ZqZci6Nn+uvxEsfp8o3LcpqBBah7WnnYDl0h
ngsUBK4sc3NG6/9DaL+1sAnqnP/BVe98ntlmxDDlcphCBRqbTrxn7fPqFvJJeKynrcqQzYgaPr0z
R+8HMOgUjae0Ks/tr2jShTBlL3DYCJo0aRlDBTeRO8uP70bEf6r3VV9AxVzuNnJwhMoF34sa2xJY
2Ozr4WgwwYk6exmCpUUEIzQHwxkmmjM+zY51wP5u4q/VhyoM+DST+ccG++f+0nwdzeA02q6ckfQx
Fb3Rj1pZWehpRRCpoBpnh5Y0Z5kDhgwUGORxNQyHsU4KKzJhkoGzCS2dfIAkqr8QiRVumUl9mL3b
VSPKPo/L334RH0JvlcufTB/gSoXJwtWptshbt1vPDW98I8zM05GZ2+Ru/GCwl1VY4QgzHIw5dFq+
2ckQTeVcHN87nIX1aORwLQ5h8fO6IJYIYl5+uVIensxNKBucMuS7KBD3ZvbVc82ANd9NQg3R28oL
BW0tdFE5vVpXhHn2SzCpQZyICWCQUN3ro2IoQQg/NDpEFX0la9Lm+5xWe39C9iW/89cJZ/xbPbqj
fnUK0koQ/NNtQ/YWMwLj3HitBuMBqREMHeBGt+IqOdETspe5AN5e5KkjN2wwBC/iROmV+t0Ze56Z
Yflf6X7e1TkYVuZl81+mlGn4Z2jcLCrWLuO2ru6AdnRiiFkV+p9ACPO+h5u1ZUNNJPDJ0YqYMqia
VSpJjSCGtwa4LXu21g/yBV665jjUMaepjXXtrVkcj4eJXx5EhR/i7AHGHTkPR8K4QBq1gCUCk7Tc
SgZhT34LOPdX2SmsTSpr9NSDwL1AViKVVs40ZQ63qQFiekkfr37J1Jv5xaFoAcwYjJ7H88/c9jU5
VmZOJvlud6GTv9b4fEaeV92XU0xTyVOGGOdZWY3E3DsAssCiK8NczSMeHKzNRZKNT9wYlURTwbNm
44rNoV3QTUIpZNm4AEyccBq/RCQGXa7igZBhKE18YLDLRjPgqCWxNs0EpOPgr2+pRYQGLWVIgOJl
hM7f7PTpJQWLruIvS3EmIOAE61P2sldM5hxU1LCWdVf30AVdFXh5dPlgKzWPgnbtpGyUIfV9S1f+
BjF03LGadD1cJcYpWSxo9FFXJYJ7me/j0UKTuhbe6NgDK3EXT/RC0Jq6t+zo+Kk995DzzqlFOBxo
xjjBVAwOU6/KUhRnx8FFtPAmx848JoWwDKV+35FV/E+TJt8OLV89kySErU+mUTUsY71aIL6Spz6m
g5e7U/iycapg05TLwGUeJJ2BmHIxGwXP7KfiThDbEzS+uN/IA5vNGUMt5hIjVsoHLHbpwO3PEGdC
9aS3VP2cDzCgF0F6POgGGTYNRb9W1noT/9wuB4bj1YCAnxM0coHhun0K2u67MJHoODC+IrthjvIx
7OxrMDjQLT2kx3rZ+xs607Y/sryOHIbGHVech5fcyPvac+C77p915CeH2usxgMw8qUfmsIF//2nI
UC+KtftPRkcCxWSw5cG25+FtFzyRX58T9NBrtd47ofUF5nBQzk4Ak/+k1i+FwdEdhjSA6VmoQhw9
gULW/DuBESBAq+Gcp3PSRcqYBU06MEVLgSxl+6RbrBxPytye9QwRGAEeTrma4I/ENa78VcJL+usC
oSwQBziIVnG1RiVUJuKRwagkM//rbN+HpOLGQeAvOGhV7/PnWpLeBp9DrEfnNR90l22BIKumfqZG
7E9bvvi88cO+VabbkvS2PRjjq7l/Zu24VWFqbHHHygv8lm4iHs3NVHGZVtg5HyJaXb6n5VcVKHeE
Xq4pSv8f24a7ca1JLhPn+HwwtGfI/UOH3ScbDPcw65X2kb71xZw3brfZEJolNiJcfS5HXQPo+1tC
uy5N2V2ewkh1IQPoPooxGcxJqVbbZIYNjZ1Pmoc/pSS3j8En/fxgcxgMrYYwLfqj/cPGydTVm+Tt
SoXDgn4lcpRq7uJypoqLO76RudJDqnuVwPpN8DNqPuqW/OBPUOjpBH4CkG3W8jKYQWjfF/QEZJSo
a6H2URzbKKtBynMCaoiwAGrplTrR5yu/WY925t5nl+DEliNaeVQexyuITkyAYJZiPzCzzzFsVr6X
mbLKmvvcjvaMIA4FLkEFh2qf+lAB1+JQHZ9qb73CUzjTgm5yEni6aMuaogwzFhipJc9dPTyY6KD7
rV6wioEezqFwwqRIzf0ygI7p+wkG/vQ/nNjhxwZfYGjrFK5+R7kuqY3qNh1dxNDceldVPswBxINF
flTC+odJjxJbkq8WUwgR5snlSiVtspKa89pJ08A6zaEUPWSciSxD90kIYwjdI/RcP4chQ29wZFLB
ZdPtUV36ukEphdKu1AJ8Pf5ZLXeG0sWZpIryTLkXSdfNgnYxusI5COyoIsclscjkDj1kEfL5c97F
jnZWHwFDczYmchFSnmSSbPk1Ig5RDq0s3pkNCyfILc6T/YMXLQ4w97mh1IgODkb+YKtA7B4yBKSO
qk4kewiUTjtrCOK41SolC253xMAAL1hQQlU+6hYRdKmSOgJn9oBISIJkynLzY7jwNvQk/N8P9vgn
4tyAPb56XwdC2Clw3nSbm5r5HCiw76V07zBleP7B3CqlWJAGPAs58Y7KzOh/eeDiHT4F/xZrHjDU
Kg/VIfIFhHZox+70wFFJmHLIBNipdHAmICqbEPbAOEXdSwMJxHTfJKdA/F+XvN/kULr5vg9cYC4R
+6WqgupX/nvk+ma5Pl6swePwm3wkDzmRlswR3QitwpRhKQ1uvYKuYMlFUHaL8H/8lUuVL1kclPQU
9yuQaYYAp+P+AqqlnDZwiODWBFgz/cCeHYYujrqdYYksHN93QGiDVVwOV1vF/9wJzi4kq1nViU0o
TzlqlsM3s+xVpmJdVZGcoANr+EhJgyOUBqgv78c15WJrM5fRCO3F6qDsiosbD2acdRDogrm5f/MV
IieMVtkz2aSlNVdcD2nPcS26wxlEqMsV1ZCrGJltKJMLSG6l7kIBD82FMVw03NpIUgMJzYpe2oPW
idbLUIVekcCOBSSS6G/z/Vcz23n6xZ2rd+yv9b8VsM5lPrj+9S7eFX9Y1EDDrORC/GysryDuPuTW
RWjvImk2vXnfTxMY7dqdeZbQDYB4qXGKccYmW9MxsUTDiH/3P1kxgsW7PSFw14NJCLwaVnVP6M0Q
ma6EotLYHqvrcaP3BlGDQ4tW0iGRoG+DDx+DIASBBLVzoES+kQzH36JNoveFsTwWEKExXPETISnk
7GKh3g98y9UsKOBshOeIKfRpL7u7zIoCjGjFQnFFjyIpZnNKRw7L1F86Yx+NDyaBj9a3IklXI/ju
FoWPrGS9qTpFcy3nQl9eGv4HfBI3rjVwVicRSPaUVLJxJcjyJ1qspq8+i1QBmjrPPJWI0gURF3iQ
vlogYgJrMAvawQFkgv70htdaqRgXuwmslz3O7tCgC2azyjJw+DShXxnw5OjnHnWFy3Ft2elA6aAh
y+nCf5qUM0v/V4QinJYScEntH5xbv5W+h3iSBKAJ/H4WsVAM0M8EABW7X0Pzp8n8jd89qWRRDq46
iKgRluepr3YHl/VchYi2Lf7Eaw6OLNcjwb2pOhjfp8dvo+oET7rYaXR4GQvgO1p/mYMhSXpAvevG
dizip2V73YoHPCycvb7B4LNkVoPVDpicsDWv+Q11vp2eunFg9Gob9BAdjLHTffIvvmxFE31D5HK0
GEtujxH0CNgSlcrxovqzHr5SmyUVExB2UaNIg8oi/vSVqu7KsSMtzdfdiGz16hSeDJi0An0rpmpO
Gdk063UmL5BSvedCaf3dVPMzsv+JuNwajCwytetyG4Me5qrG4SSBPWzAyfmnwKaRu3qJ4XKzCJTb
Qgl8tLmf1oM79FV59wVu+CroTK3zzss6duUBLEWLZTpUb6gfu0QX5JqtIJ6DxwaqqUOQllSANRTf
6YJXSoaaf3cxj2R/9h6vw9rx8apEzbYAedgukY22vbfrQHmb5G1UUuWrJ+ctU9WAl8+wi91I7y2H
s+8AxKYpfGVoAEaVPiJZl0nuyOWlvbOrXGOxXfT9g6V2jqlfWrZf/SxLBXhkUpc6Y1PUbEbdfket
OwnLHYG5Kmuf6i1ro6CINTh02EQv6ku7NpxPA9fOu6dOZ7wVIXCQhO4XKxiC9XAeK18TjfVSA+Y8
cZhVclmTDBO6tfPsgQHfB5TNID6Hdo7rfGJdy+x7sQXPiHTgiEiR85M8ONCYveHKhWUxpoZ2RBGH
5Zlj+6GpHcyvXHdJ2x7JL74rH5cX+14YuV75LE0g8C7qjMimHzzZDFc9d5bjEOHyhmW2P6kkuhOf
vlDsV2ld3MmRiVKWgSlFP8nXGGsczpscpcwucavxKIm8XyeqetBnrdUtPipW9UhkE26DuOIVh/em
//U9s/cBhTE56XmGNgcK3TRuiMcNMJ0OwKxlBuk20p3SX34Wc62ux/+N0RF4fEGa1nTXBqWg/P1j
O8/8Pf+j6D5YDTZs0pQj3AGvzJkkqJWhCTO5X4B8yZGcr1lzPaeMF+HKC/eFKFr+DkCD7oIFRzjK
kYkittWxye2u2U7SpEOn9DELn0cDxgc9zeDrZYRkCa4hLfURDy5cH5QjX880sTkdlRDITEdUymLK
U2y9QWQ5rzl2k9v8E+w+2V7QaKfEKaLAGKUOBaEw/aA+Z0gQxHlOVBGPKJTkhTQcRg89UmpAemrQ
b03ZIEUZiNEybwjb1wI3ayiN8BrvnWHFg0oMXJD+gvA1h/cw3I1w4A2PTgNHfzbVCJwMKHxdIl94
PkBKLikRCzRNfWrUo1sLW62A2VhA5KgrflUbI6lM/fYRVV4Av+Mo7VFar8Zh5dhMpeuVQ+1GmS2M
t/oFWE2igfza/Xp1MhEGPxoWK+gYQEejY3bGj5+3EF1kg9gzgx/KMmRBnGUWHyMpf/gB5vsWRi0T
itjk1SyTVuR9KL3vMjcK3dOHWBHWysdn713/8bJeD0MDZnZhLwx58+slA3tt5aDMkodFLwgb7BSD
W8hb0dKDlWMKq+Vqh7gm/W+e5urSxuyrFwcEd4GZfmKNY+MBPRqufx8sjCTA1s6ySmgOlkBvicrO
tZ4cw1y9Kyo8sUnshrvDGMl4y2afyPQCcKUKTGGYVwAUogf66hMZ3OClWWnFfDiuhxm1yayyPw45
GwnewWkv9pfKp1jZdywYr1oy01ILEy/AdEh/+bFHQwKbTQclazaQ45rEgbszfUk3cVIz75R0C4pk
fhCh8wXZQ1WnUYRyixglIACe17GJ6Mj7bEw3ThZ0JOWa7xvn+H5x9U97LJie+82Q0bsEmQs2O1yb
Tb6V2eX8a5UsBt/s3SPxsSn3Za8yYI4xHbqAqAXMWiVAkbT1j/F1qr8I2ObLKUvQrKT1jhnXVk4G
O0nw92/h/GnXrzwbL94Pv9guzRP5ckGJRvav0guzRI2zpPPebS9mMRQJMMQVpbaU9q6tAs52ODZq
eVGsyyFfUMCys0O7Fg1lDQsXrMhjsKWdnLJ0HkFfzhlHFy454qLAJv3rB5HvVSGme2AJxE97f2l8
2qLa1LMgGkd+JEHiOE5MUrN0BRHrLceVZYa5gYxNDQfpMfZjYBymcqPbL1iq5d+Psx2FGGt7EwER
9gU2jntTbBWjX5H6PTT0ZNOxoznzDIUeBN/2jyKpD+gZ7DShq1ZG1wcbM4XIUpGe3czj9oDQqoOs
QTxBsgDxMM2cZYfgPuNGCoW3ZFuD3fdpY5YYDy4YJ0RbVYOuBc72JKgsgDQ2CdmN4cg7WsAz/RRy
dcDgAlh7FnUGrbJDhVbNZXwXkULCz4TKJfLnkCivauNmmZcrT0N7Lym7++Wg6e+jmypD/CJw3PfA
E7OztoK4psm/3BFLxvTI5ETJV4Y8adIfv16AfRowTRK/EPZkv16OFeY9CJfASF/TZEcfrfS2RHAc
9VOGIz5wHdFTTZH+z4Cz4kayeLwo15BXka+jlNJ00VvA+pG3QbCmIJZb2ARguVr/OHQus7D/FwNN
GPvfIDYsQlGQbkba/udZsIfAIEvC3EVECMEf6C6A1pT3JyHkODVBc9Lom/s2ytFeNeM8qArSBEDb
zQQO2UNHRX8R57nHRcdcz4zdsTxYAyLArNFmh68tuB82CC5LubZWXeXCgOVoS22xZX0bm0KFg+cs
KUAr/Mtt2eo6yNPLqZj0DZMbDEXAqf96Cm4CliAZogWnVek+pUHAxqk7JR/ysdSkSuJJby3f7Z05
i9vfI8/NHOQUDKLCSUb3un0JihSYQLzJQaIs58mYnNe7dvEVxN5XtJMwVBnBKlu999Qz62G8Yo7v
U0a6lZu39SoDEm9QykmCjlovTK0HD73LmknU148I0eAGNo+m0y6JMdNvRCGizvR7lDtSM5/cl7cB
wZeHoyMbb6ZdfPVQKWqOS7ViHK8X4awf9Qz7OeKCGuXFEYCklLyOcHd5ZU0aDuzB8CSkEGwcYT2d
qEEu/Gp+j8rmPAtNET4WDzDzGos7C0dO2Mf7mi5IEuyQNtMKB2QdIMiltZEeSrm8aibpMIND2Ot/
Wgyk+9KvkjZCOsbVOmZ/BwMAHb2lnngBdfCbyqN3LbN+hj5O23GPSqyPJrWjQW0lfxlZhC1OpCTu
zl2SJ6wk4y983Y5BD+XbnGpMCZaCvBltznZUA3O96ZLYhBLvarmjn0ZP0s1P+P7AETSXqtozEOFJ
ccupPTJvam1XeqvJ6h6ivNxW7+0t4Nm9FmiJXqIEXOXeHmcBWGzfhqOGovQ1264VVymr1LERPuEu
0yIGIRnwL5iXSlQBeOzJ6KUqpXu5PqtYtIivuEOPtWUWZrys6iBZbMxC6NFDgTlH8ghwEkNR7AKe
0pXS4FhPny/qZgQXEwG5Uk+kebiwx3LFzGfEePig9oV4nvNhRvT0XbsE9ZbbXN+sdlDxkcbXD2pk
lxc9nGo+YiOaZqHhpDbwRhEmGSdxjocS/H8/IECK0nHO0GAsMKxSKfbY9z4czVPrbr9I8xnFUeE1
jUYg7v/Uv8T80aJqeIBmLnfHMrezeIrPMt/MWokUPVrX12Mu+jmIdJwtWcmyjXE1RfLTiYm8d9CA
2V8LEUtGkYC+/q/y0EOwiB4wvQzDoImCc/axjF4VEHln84U2T6p7t3B8dAOReXa5TLI0O3p4kwiv
P+xOGZFkaZ/a43uLDsxYuWkp8mYWjhOWbR06McYd4ozxa69tdII8SGy7Anl4G64NH8qZnUMxL1Eu
p7rdPKEC+IJasUxfOR8eDDwWRH2vpf1riuEPhWEswUH6A6qadcMMWAZDIUZ9ZAYl7Swul5S6LTOP
wNiz/cyo+xVWbCz/LKkXh3CX8/pyLW102e7s+QtfX9ONFOs7oqzW+WmKUtt7gOk1T6IlrFn8hdxK
6R/BK6hCVOGseEkVv5CrvT6hegh3GXVyasAwitW8mXL2bkUVOaUGrvbb17HirASNwLAjICNJnjMB
IMpzcoK+NqF5q3dJ9eQNL/cC6fP/JYC34daeh8tu6WpxH+EoibrC2DGvg3RIkrnKGjDODDgFhzyQ
biCmgGrfZlU7hLkP0SwczLtCiqyAv+Ak8y8xh9J9QfyELKEm/TVp5aH2bH0k8jN81U1pWixDR9bu
62Hi0FpNdgZi9To2HPLU32a8wIi05zuk+3Ee3JPi6WrkgVO3qxFTNmaIVWTihrgH++ebLgD7tqG0
o0edOdo2oxbrPoni2Gg4KS44am+/Buc2J0q0YnHuDkvXLIJM53iDm6DwO+4xanL7GjzRduktvp4S
5QD7aYiYJV5HklPYeeDjwc9UcydJxXHNx2FKt0dby0BEzDXbJRqg2RdA2wH7Ox3jyGQzJfAfSQqM
iGqkfDRpoS+y9mBCww3ZBg1WwJ0tOiXNM9qzAvb332pu/9ZidwNcICblIIQ2hD6dUMjC6Smj5+5H
IjphA7zgD1+0+byzTnt65GoDQAQ5eqOULtiLea55G0XA74Hgax7yeyUf4S4j0bX3fXhdTr5y1W+W
bFUSTJwGqk7lwZFma0nbqmoE/784AbB7f/2+xrYIGDqvMa7V4NuwYxzu4AARkiIhoTDFw4YRNvqE
rT8a3uP+2cxUXEfFfA2YPB5qFnuJ3xynvIvSmLrv8Ssak82A5fUxCI/lGzZntgVlZAE0kW4zVfUI
hIwwBj7b8Z7JXGevbl3Z81kcPU3JQYbOym+ZU2Wd3CmEKwgySdVdDTLo9auOA0MTAdnMYGoguzps
DT4iBDXK/+4blpaZrKQHHcWKaITL5qDcEdy3J+RTpHBPq4fYPX5be6KBTPdxLMOZxE1IfF3uz9F4
XOhFRYQMM/7nsF3AWDX63Z7ztgGlyTnah+/EWq0LC2T0KTDaQWaxA3+pm2NbNwp3EADaVkSuvNFd
s1/cPf/pb6Z80bByp7GyDRiCPzHi1FywSkAx8m5DsQfhsuBfpf1t9+cw42WOf3gomN9kDTMmEFFM
QdLCPmcqZXQCttUBMERmAWf3vdOowAAFyEqGNiBGQOD2zF8cfACDhdC8TAmTMPjFyUf5D9eOo91T
aDmYnl5CcAy/HQRUfndoRLXw4TkakcwRL4ZtJ0Ua8T4wXzONyBYX8Fz1GKshFQsSbR34cXVzsVLY
VY+OPrW6I65IxIEE95V5cvINr/2h9zJNoH0Cf3lnhv8JsO8IvJj62EhRlcoXvJ0rizVl17ibmkTl
LZLz18s8QmKmnFDjlxLZd8fPRtfpU2NQOXzdkiq718HNWfUj3Zr9DOMgPNE8BjC0rXKYDr5zqkjM
jYarfxIa2Xp3NEMkMUvyau7sxI6BMNqakxMUmddE/UEUoJDwgYPWcLqmWbbFV3dSKJ9UU+uMEk7c
IwJ+OxWuUUO/hXIWnKESjdfyBLz2Syh2aCwaavE17vOAr/WZEfly4ugVDfPoDXw4utL39Aj94EYU
ipHnoAz3aUe/WUQI6ea8cRGzsY3d76Y+y7YHcGvKWoBmUnUX/WNpKtPNzcrGDHgSJeiZQK3BLdbe
tNPIU19ZEXPbfporcdS80c2NBY3nQGF0q+lAj/BmCSsA+D7Ff9H/9gLeaPA40RfW2+ctIr7k8Tiu
pRAROEfBbpol/FDQLgaQR7wzkUuPzaWLSpZYgDvfejURUoMhqyxjWzoGaSynddECrm1vvag+AjXZ
WvESVLgMjR3swtm/EcVYCTGGmTyUF1HaBxULwS4rHcyZkca1qGIVUnYNOqDdxmbRqUZJi4nHIdkj
02BDi4m1ZoUFGcE/8J2loMs/URWTtdLc74hjwpTw/OV4oPk2OBRdNM3RH8O5v31sl19f8YbxJ2Ih
Bu+ti1XTxOowo9mQndcfhtlnmQz2usk8oI39vVi8m1x6OvG2w5ScdZGMbDUr7zS9CwAILhYuVlWk
MQtZm+52yffGhlgs33L9pd87FDjUhjfRNvyTq7basEqhhJlFHIHGWvJUXfR3t62eZve5U/v4sWpI
ztlD8COh84/yZozoTSk+XzuMyBmgx0LY8klWdLoYdoJSIA/W2xvdLjzP4JFgGzkVRLkXsr+JLuQt
ZC8Xs89ZxND29Q3e7zz4fcibFTRtGqmTWr77Pdd/q9KvSrHRXBwGTWjVjvazrx3u6ih/ftEaW82G
Sr2kx6QzjdqaPNFuI4TxZS5b3I+CrOEAQ43PcNLZ6N+xsIF+ISss0gTWsSpg33uOVuA0BKmFaezG
bjYLNF0F+UO+w7SOaHqYqkZf2UGWAE+cuGtMTnVAI2Jv8Dto/Lqvg0XblqFhefiiN39SslNilasD
bmpuqMMu5urbs0XxIOIePbcS0x9ai5MYn8ln/U793AXoHlybBl7NZqvMOx59Cu2qvKtOLrLOCBE5
FdBFaOdcC7MXoI9hReOHRcauA2GDXEbzVlWBzgnjq5kLOLkM4d+jQnxuBMXn2eFwUKSqLga3cQG2
L/VDPX7bsh6mDLMPB1s4nEmSg3Ps5oTM3n/vfSXceBFbJQvHYhC5ZCQtQMUoNMUH+zutOa9o6vAu
Prxjndg4s0pX2BTChKqTKh/YArepL7AhqDeRm0hEoIShZgNLcd8wWfRJFjSggaa/0Q1ITf0uD0ap
FCJ03E9zW6wrnd9vp0WP4F/+cGk1X6rfgUOLcfzi+PmXWw58uP3bQ4huafzsU6LtWttRxvU+r57/
j5GaLYtXn3OHmw38GWWJIKc8iOxpxSh+qD1clNv8v3eeKRmgquVVh/qtcjvZv4G7fcaoGdQhGo7S
+onERkilmBmDa5wSFnHMqHKQoVgXPFjZUkTCxOk0tRXklMHmzgYAeXTNGCKC6Ve2kcDbBtbD7l/5
Nwq8xJIM6ln+sJ4QTunMAd3SBtk7kTmgklfML6KpMdyp0/1vlxWLtghyrfRFgXUpIaHS9HS2SXep
OiANydYlfqOGT/bUFnSYgnl4qlsPzSqVccxGgcDEuubnRVIP37apYK4ACF1RGjW8Ynj5v7h/2+e5
QSsC91oEleYnkSonmzOn+JVL716WYCewRfsLZlky+BZezm/A4Iy/Vcxl6srJBFGXD8us7/FtjlH7
zrAtdWtAMfzFVxt5A5dIgso1Unbi17hazwEF4Z+oSRt0giSv6tBSyAP7wi+p8caifpzLZBis6W6g
SsPFgLZmKKenAkmb0cKsuY9H8bSeOR5AYdmWp2Q2Oo/Vk9ytWJNjViQMqxkjvl2QYPAUYiNWcE/z
maw7YTRJ2lSrLAH10Aodz2gKt1gT260sYAEk4NMvJE+BjV07z0IBwWS5XoQp0pHZF9gMpJCGfrNE
pdXpmSUxOtjKhXgYnB2CmXPpF1HDgGQIDNabcumK3Q/AFQwB7g536SQNqdnMcN/F+tdvJIP+oleV
HjmcYlwyLtYTb8Id9IF4QK9/B5hWEE8WjOlMQCQB82YFYtaiwgyUvKRBs4X+pyQmnLzHcdaI8dh4
kQDQvwrAar2AFJMzxiBbhjFRFewmfsiZjsLHMys/As0a5zM9r/3++Am1hj8PUOWwDW6md5nL0pnm
fiHHFFaXxfN/rikdjGZigGK++6zjlFKJI/gk0NyS8AOidHVxhU6h92S8ZAJ67SfziVvEYdVLBxMJ
7MDDUXMgO5u5GaNt0nmIildkkVx3NxA2+VGM4c0GLFR+FoKb3TSoR4Ns3tqX9NUL9JmRkHgeCzvK
RPMZNJykJnNWXJ2M9i/X2cIM6L6AYma4CWiTNDT86lGYN/TlJtyCd0ORlTqmPJNkOUGlL8JmdavE
oVM6NoP2lE19FPz8bc49Q9iWcnejHWs4pNvGOJAWxSLhbJyV/rh8LUc4pk4zqsJ1Q3J6K1JSNiKw
qMqfDGci0YlQow54IUQFxYVC6lWPGzcrpQWE4f/aEWqkaeaAgH/nmUHqkgjtGh0uGNkNdmSIEHmo
CZ1rfxa2wfBZHu/MyPOmRwEkhVv33Ewfud8hlr4ATNU2wlwr7jGZpwVvuWzVKILHHX1toSPDyqQm
mwCvYSbAHPgt5xJf7j7u/DFszDU64AgYappqISNwfEg+OIOV8i1/KWzEHUe4EWxUrMUBEAIPFZXR
ySxcN8wCzq+eGSRoI8qEIGqgdLuQsTe5vIco5lZAhVfJMRnZuoi8JRFpsmxsPSUQ65obPBHSnB6u
95umRONdm0bjTbVkVFUjKMCGXRV/sE4znx0wPYJU0RafC00NxwfprDGexBw42AgoIuZWisBl+WcG
lSGAOzFQExumUsOWeVbHcv+ZYc0GAdmpUB5eSlQpIFbITkOyT5qUNGFh8qDolA3h4EGovFatE3Sv
e52tfRYVlZTu70Hzss+Hz0QL+br+NtNoidXS0I5gN+OKr/UcmKKv9wMIh1iOiHn13RnhMSahzrLi
rJvuLZsM2PHvfK6vzfxANLCODNZKVRGK/rQq/YHVaKKVsRRZI67bI473c3/clA5v14vCcYrvtccC
ux6SWZofZiC5Y5d9sVyhwKKyrGTPjNGa1YR/lM1pEpmdAeCToIfCjeQi5QEDEheEP1SGs4jfZhO6
Xxswak2iQWBs5jam+LeqsSDv9vwMr25JMR4aSfOI8zalpxvlMfTvQeN/5Zd3JHeq/Ciak9bmkOFJ
5okd9toHdJ6iQJmDog/tyKeR5JDcFHl3fSJNp0ke12SHoX6Hswter7r6TNuw42Z01bLETn45ReWu
W3umJkXDI4a3RrXJFbTkJOr3tW0Wz4w65Ecsq3oDPH15YWL4LLTgxyDppaE2yT691RbNwlLckOoZ
zOIDrQDyQEgBK+nhO6/lO5PraemxD56JXxgYWxgHVpmd0s+46z8TEmZxQpnh0lPyO6Rm+EJtooDq
6ZoR7dyP2911Ucewsyt9QXAzB+eoFbF+3KwIiGbyHYqEMSpbmljOmvpJemZwnu5qq5rBSjWPxyRh
a18AqjKQrzMzb3OzlXFRvxaMwME/qxkhF2MGpbVNog3I59OlqO71PMQUCDuOkRT/D4grbMcYCzCO
w4FBfaVXWGj/kDAEWhWeXHf7kgIUc1rWjPLz+hpAr8LWUcP9CRNyWkSjG/JWnoiMqjO24jjzeEga
wbo4ya8JBTWBHyBHqIHKwkPApT/XKBnQXuA7GC0/pdDNEJgtz74Oh9ebddag87+/DczX/72cV3uO
kc2V3BKPjn8Zw+ylYzVWdIzRi4ETor3S21sR84DHrI9Lw5XYa5cn11e/30cZqDDKGdc/JXFPTGFa
axxlFaYqtbuxH+zntYP6PNnHLVjbLmigN+0JSO69yZksj3PCnyyohZMxJyKqxAiPEOoErvmgF6yP
NBoM9PZF2C91wfpJJEFUuqLfzx3TaFP+mG5gcW4jTjgxa+tomQ9ZG76yKuFrDWuYXIhqDip7CYTs
LUkaOB2qzt+2JXlEq+dhMb9OvQdzsOWLMqpbWKcp09qhXwN9wgoJqG4MI10bfLeCieKL0Quu5TnL
R1iKyluy+OGADSLo0cTTuJwVBrd3BobqNruzUo2f3RcuH0PT9skpECQSkR3T8L7tSO/4Ov6q/mYX
yNU37C9+Mc3ZY71XPz7sD8in3kb3HQl5w2FTRd5tR/3MyoTIHIjO/MnlsSGI2qcuB3xienfV+wsO
W0XGYOqh4v9rTtIpvXQfRAjgqHKBmbWhOSjSNvV9HGvE9/WvvL/zNrTO3QHIoxpBKQEEnb86NUry
vUAU4RR6X32y8uhlRRhxMwUbZo87lKrFQMTxuriW0BNSo2hu3nFsjYTLY0sZi9axMp45brgYWy0i
2vHtyzAHdakcR6RgorGgwTWiVRQfx3JDArdQLTvuNhdoltD4eKE2+bw2epag/Clf5a9nHhqKFbXr
cZOcmNjS3vwvokI00sasVSdCmlY5L6HyVjFfdPKxX2H3G4AGPtfrvM9/bd8e08ArR53SpH4YXeE0
+yTPhq38/Hizbm+rb07XwmHbBmqyb8rWrcHPHGxkRLuF/l9OXC4FLNVeJ+gBmP0zXiFY30/SRiRE
wYevgvxb6shDoDkwPWaDbhDukQijwM9/U8p1WaPWdHsx4CPz+roN6mkEAuAsY3MyZXmtXnGHJMhY
yOZ1O6E5SFaLQL7LKiOJY19i0o6mPwHypsLqdU4IuMc6/fNpbtADNt5p/ZgcC2mI1zeHkSy42xWm
P1jQIoZ9RM6NJCt8xqe3zR4HgbehPsMM5j3tL1fy0gb8a4kBtH+fgcOfE1HPsapcnhtv2/gQNxF6
vlBwmDOFSXAUw+X8P5kwcVDIE+GdfPWLaKpuJQhyUhjy2o1CcK9cMIDAT3tH7814IAWwylLpBfKv
mbTlXEbk27xvnElwdRJztpYyKFzQ2ZEzDZCuNiQokmPJeKLPJLUCRzcDsZ2Ym/JLrU8XieYl6s51
i+3j/TfQrBDN81dV+l5jsruugDABPJOICACLL7DI1v22Y30pjcYsfHdQPFncbN8/c1Z5PEFPSYU9
fV9VrZ3MHlvwyo1PJ/GboB8dys7eDsLlYg8Q+FWUaOoVPbY+1MWoWydkCcc+Ip6B4c2t1GNyKNX/
R+FRpqa1uhb+Qstqnrjh/llMrWkJS8d3sx9PsIbOB0zpsO8V3oJNtZkYepgZKxrAiUH0qKptQ6SK
u7ZtB5r9MckMfFZ7OfNFYmNF6+uV7qTTPsou9/yB47pK+JD2+SwTvaFaySP68DRSJrA0lwFbgL1Z
Z7YtNHjdlmQ3iuzASRfDxK1w+yEbh0U4xGtXbWuC8hLqwOMQ+ko17iTY6hZ+aLS3Abjprfj2I3/S
mwcEpJXufxL3eYZW9KIsZg2RYC3xg3wo/MISEEQEgIsfJ8DiCnN270fduY69eWTB/BbpRIyRXwPC
BwwI6vv5Bg4DRZqsMA6aCTnyn213ZTWdFdKO+dO/EKUW6qUslq82pValKVRIAyFRdxW1B1EGwNmr
wjiS4xVlJgg1aayZfc5D9NlgF8jtOhtKjOAQ86Mgyyok6fBF2nvLS0dwBmDg91JiH+OxwewIleh0
2BoGVOdJAYEmv+4Ob2/gJnyPwtsovp6G9KKm5XFDYcVBfi0TZInr7A3jDZce43bvmf3p3VFFL79c
quPss0AyqZ0kt+spPKEgm/sMqWOG0jDmYtyKqpmZOgxz2ofr+dUtHXqfRb9893tDLlq6h41rD8EZ
f0iLZ17nqiwmsdQ5IglT+8WgUc9z8Zkthf9RVo71v4CI9sLgY8Q7zh/XE1WfuxqctOrGU5EeqRls
iys6jp4sBKsD9ww5AfW2vd+78IZqYWFcWVfCRqu81tPF48dRerU4B9ESKEGA1DahYFGuIaOBTOD1
fC+9A2z6hRq+qHaaLmIG8N/Oi5gLHpZIPtt8nVpkeqKzLQ3pXcofPdKapklHlmknCLQzLsuN0YCh
zwy4pFiu5A1DIs/c23Vfx8t9X+Wddkuk9+pMMp04+NLJAdGbT4eF1MzhjtuLIEtmoAYG/FN5DJdq
UjZVIsN4EL3OCqljZ2zIDz6o1gSeXL4pTSCAo8KeZYiwCVmJ/7bSeIDgUM9X8sF5cBm/Ywvu04FK
b2LLtjw6fLFNCy30XRZRonzMsgQT7V+bIROZHIQAmdlehJWQu1hR+9mKDtSqMHJV67RGEE6obyVF
3S0Xkn7ZgR8YV9cqfKXzcBH63lpCfvKs2S8x8Eq9ep3ERfh7EZJEk8Z1/nMWyF/cIidNiiVog1r+
1Jz8LajRE69jnsnDi51w13lI/R6iDIbGSuBLK7mjMQvzaJxidMD6IBJJ1Dd21srjdg11X2DaDIPl
KIqGoV/qjHwMzOTErx8QDjbJsSJDo0+2/opuFw/bjbvkVY3A+JVnneWAAMkAVixqxXHFmT+hX3SR
+h3FNmYptI5jf6QtHkHNAm34rOHXMCY8PJX/vhUPaphtOsM5P+DijMNoqpteRssJZ3pxXCQiCmYn
NompimtF84VsEkCz4NRDJH2h1lajrganOb8j3hgeKZXK6DQtABvW9edTW8a/qLTPOaGwSk1r2Prc
qmMVWpQo0uZFIimEyUmGFBchL5t/D48kDoX1SjWxCYnqhBA96bd12h3BfmR+7tLDAM1EvbDWd6kx
L/MbXxZy0DJOk7MvjbaKsAYi2HAYp89j+qjYXce70PJOnDka+VBcsTeeZzQUvk1dNfQyH2g/K1ET
GPmJ00y3I7QRnRGFe7kiMYd2S+CDHS4aZZD0E6wjE2qTn4GO//oy+8Xw9O2hXfU3OH0Vf/xkKeMu
bh+jGyIs8zAIgtC/+/qHsABiTZOyAglRkKWD/dUoCOlj3nOwvZEvcPgjbnup4RaFZPzgJOvnylmW
mJa9XIyhnvJStBraBjq3LpvK6vkQ3FvtKBNMcoXJwYxpIkIWzj62oaDkYqrthqCgIrEscpFxZIgf
9SuJZikfF1C3e4q9M5cTPfahU6GEQeq9NeUMm6aQ7YOOc96yfKqelE1nuhDbjfrxUibOlzuc2KWW
eNjYLGJlXh57gibUWm81O6+tjYyXGWyD/9EU1NVFMJU368Hf19iyH1sVLjVORQRkbXuFzKLoh5j2
RGrzx3zZmFod7tj0cvgln8wI9Do/0J6tnqZDr1BoXq0vsgtdTNrDQRrxXIYb0241TL5hjZqCcY0a
/rr53t6ggsx5bYQJSYQj8p7F3EAn2BdDjzXBEIh3ntTM2ite6fhZzg7rmxDmZmUkNplFAe1rMhIn
6qsc/UvAl9+xa1vxIhbYGoaXJlEhxdAtEtHQ+8rBaiQQ9kbijS4qYxwhYjjv037EQsusI0MW2tJ8
rZhJ2p/GxNvVcRnLZWhHkrVE6Qwf0uHPMSQw1cwWTSOh7yELi2kmPIz7kHUiHHkB4C/aOEKpTlrm
sHgm/V2NRwBO1sgzjDZco6iuC0waKoiujksvtcaDUzZjns/L4YBkFARX7Q0uF8RJAwGSyAni6YW9
PwjfbmQ4Oenll/L2fojdvoRz3/fbizaKnBlx/uzTf2nekWx3H1ZY1Tlom3PHYCmlZAZDlz3knkDW
UbJVPeFacR3MYPTsYw0jAMfHLiTcqnKd8LwQEhKCGga5sdHTowtgntmwfoPCQuVAKvAIVTapbcvN
uw0I84vKSNVpm3QibZ/lzCPnIMACq0ALOk/ng/yxS+Eyrw8UlRxbrAl9ztbOvLI4smqp8U4imaeu
bbzQfyD2lGN40IBnByvNy4e2GXjI6+edemxuhqdUI1c5wx8GSjFt9IehwLWP1BgUOefHUgsftFUy
vn2qd5LtZMqLi5T+DYdOmNetw12ejejOMS+QzaaPeZh723XDpdMYVqA8ystTs5cE3ax2jGbkCgYv
9sjMy127tbgJ+oc1/KpRBBl9omL7YYTXoia/ztiTKkRn8qxdbMBLYe3Fh1PZE/9j74OCGzaNvC2x
e4tGd0L2m8i8ZMi95C6+IOjUOpGmmw4uM0f0HXmD9dQrvzJ9enhqE4UQbMwf53It3IpnaCDLHKdH
aUTvVvbprX1GzfXD37Hm6Lk1pEW4yhl6+GF2Z++lkfx0qj5YCxJ/gGX7PBwxCUsmUrN2DD1ije0E
kBKPJTKeiRhmAszhxVBSMOeqsLiQt6RbtE3HaoPrRwcLBiaWxvzw6QjVD4j86a72cywyBQ5YJBoh
uJj72kCA0r8hQV2JAVj3TRsViZbhyX6fO0qjHmYBSFe4S32wlVgZkBBfRKBHlVUXCAHynfecF+Z7
gnhvOQIuzVsSNxD6GSMTUg4HYSGHtV+nNCfEKFu58xM1y7MH8lVpdLBKj6T5gcLHJL10lZx0Vd7/
oNiOhuBIAcnzaWIberABj7FaHKhpMrpRiKzpg8Usf/ikfBT6XJWl8DJcQsHVpxklGrJGloLXRzx4
t4qcp65OfH0uopu4cf8ZSjQ519U8fGXRTPl0fOTHOW2vCAxrLftNdOl7h/BFAlXIRVa+5/TtHeNJ
rDm8J7ryNSU5xkghnMkuWGy49AJYrvrsY/UM5d/fwKLYLylmXjOPrc4e559naAHvl39GeBy2wpoL
Wt8bhviwlAtS+PfrDQPxF+sc8TDQVSJ6x/4cgQHoqexZFaUY9p9orFQ3Q9OikgIEWm5VjwgdoqkN
//1A6T6QIBH27NcXgYb4553DLpcLoYMTbZ4nC9CHvBbJVl/PbC2P0SK98BDKwQcSff4zF5jyDbwb
h/NVuXNdRSf53NVScgQGhcS+S9ESZHcIt4gpdnVDdpG7EB22H8jJvSa5d8LW4shcloHZkJSXGQNu
Hk4olYHwBo2TEFXf2zCcq3kxtZBVfDGo3MvMJQ3xiUL7wDUBGm/khcE8to5otcwb1Xsfn8OlEID/
mwrdlv1heTCHynTt0wVeDgEhvnuknZiEFVNqx4S+oStp05svLQyf6ptWn1ySFunTVGLU1lTNSouk
T8x2COATzycidbpQoDRIRW3SeMxdwBUZqvs5GEQvlXMW7MJ9AcpS8YLR29UlfN190BLNJxxicW9y
sU7vKdaWO3RXxtKIFLV6jIBBRV+1NHZefw2mW/dzDyaGiIw9UekmepKFIRMHq39z/4mFMXGU4gei
LCOYyL6LwVzjV6QkzAWDN0uBgzNuGKVUUuf/E3hFrCrZL35NjtN/pommaONwjsC6/VpWnTEL7vJl
augDiq+ADGteSEu5I3efoH8ouzb1GaB5psMQfz20shwVGC7KWIhBCqzxhYeSINpztj/bEuXhyARG
tWVPzkbvvKkIwqnayjLCo4EbHtgyzWcXLM8YA2fJhs1fuw611LV7zY1zF1UjtwKM/fVvj+jjKFVI
f3TXDntEN0kPAJxDJErvdhDUfJLVup9YyEtCxQPHifGU9uLFW/ElY5c7OWpO5Q4rJVJ7IZ1ecfWl
T9D/neqQlcEZtsN2dmnzhjasOeNlRX3kmiWWX880vZE3CZmGNli9VklP0Wit8r62erWHDvmkrQrS
48Vi/LLr2oSGlDkFPZrqn+qhQO2DGX/N3XOgcSDYtq/Ekah78/nOfQ/cVWbveu+WLSLKaSFK1xZc
ILg05QCQpmG2XZ+rzW6lHLNa7IUMwX0PNnYsmVpD3c8GfhL+qZt7uOrygBMGhR09thvh6zgZSOoq
2/V/RQ25bN2/McSVfQvSi5sQwfP2sGQ0lu1t4MQBktEZ8aeqDZbsoa7evjs79+k+PBnhxc3KkeNQ
6cKVakY9EGtmbXdDrK5PgxRyMnQ1EZqvCsd3YE1TJ9WgAk7lgEggxvdmg/MDWAwq2vgFkEMw7c/d
rKlUioPBWN5+dHWiZhR53SnG88dnp1wVr9BEsbf2aRd/1Lfi1BPbEiht1tXTgK0CkETK4/Y9aoql
QaV7bHfcM5LEDslSbzZMTMgiVU56woQYGoAX+z9GNy80SJLXxyMmoDrOgZdU19YaBRbIsxICHoJt
C0EE9JpQ7M6cgAro8PIXVO71S8k46swbs2Gw8w4BS4puYwYfr4YMwScTLax10Kb6PA22H+pCoVoi
q6UaBfF+XfmIoHOdiKDmVGtFqAT2SaZ3eR9BGXc2R2mFuT8+yxumMu4tTHOidVAVe7Nz/AmC1s3s
GEv1t6/92Ax28+BynTE8MNbcyCzAyXq+RRFSkq2vl5PiqGGBC/xkEFwxjRZujGuND/RPCS0A/zub
GZov5NwrlkJsvQGd6r6UVRSHQfzBuI1HvmnNJHPwWNDFk8kVODwyBBkdOgG+K+/7GEQUEaN15i0U
ltsOFySp8dLI+Y/48xdc1ndlbJ/rZxewMMxh8q8KoOnwcojwLfJnJNTAQHxvX+sQNK5I0Ge42o2z
OizIWkIW4wQVeAjwlZK1vFrfSeZL6OjXcVkMUs5h8yRnOVWpXqzVhCPYcMzMtBZrAZ+Tyu8qSu37
dAhEM7w7UmYZZ1jsKmydB43QrahH9SnhGzm4btfnUBQQBw6UpXNKo59qI+oPPsL96UvCH4DJwSQu
fb2nKMiwujcX+TWTzz6bo5xumwjjCNb1ShfUTR/oBiqaSHJO9oL6Wb98znIvoIY88S8S715rC+Sc
hQ2rvSGBAXDeOxUouNTzm51kT22ZOMKXyD2WNMBDW28qDS69cuM6vzsLArXHppaLylR2mCy1go4q
mVCbfJnbSFNQ0r4PtD+I33M3TpYDqNEYVjQdSEFUVea+M68O7lf0sr+W1CD5ZYVPpEFycCSLyXbd
E+cV7Y13r6RmbT/jbFtWffbe0bnUiG+EJf4OQ1taMH3v+Gb0HdNz99lOWNLu7HW7hqhPwO6uR9b/
vnbiZo5ovm9hEPekcCGnFL/88FDGeFM+DNliM3m9zUA5wFdjM+CcArYj3j4grg5J/adFvaG3ZqyW
qcDBcxYtSkgtTus4hMqPblLI0MdhHfTBYHCEZbhSpCCsF/5KTL89qS3JnNkXtPwS+G5Ipkaq/9gL
rdmg7x9zNKpJwBDR1z7HaDNcv/+FfoMzUCyTU3cCHB1WwHFH9E0xFtcnJKIi99/IzozWxiHUgLrP
lRGXDHw7b8ef7EYQACq3KqgvFECwNS6A2aEBmQ7iWjYpYuO+Ty7iRA/g8x1cHBoVmV9Hbxd3oHV9
zfMsfClfBcylhLHo0oeRAMYeb8m51Dj4ZrdyCwAmHygLdVPtZ0QfVgNJYJ4p9lib60YBZUy6ZSVf
YxG2iLAOGZ9pMA1asOwuwzEt+qLYoqHwp/VEvPKimqQTRVVimeZYV7wREby5hFIDKNgLi81t4X2a
of0KdwX8s9+BUu4xnb7mNNKVpKjNYytXjm5wpA0zRbMpn73YdTvpmK0Im1Xi7cgfGByMosddPwen
fFhTXWMXYCXKgO254xN4UI1qJb2VM7xmziNsGSxcqY/+u59kBW+0uATJjvaQ9cmYLcI9/YUgFCUY
+0dwKB+YVg+kb/bXiCCz/cxsfjOuPRUSwIx3ezWVVHnmKbxb5BL4RbdmNTAaT9prHhPpt3iPytSd
b5v4M/rzCPtrQuQIG/8Q485qsWg0yuPPXAH7MgQ4wK1ebT84omcnoUTaRNhp1RvZ+iT67p1WEPfS
MLv5gM78/ikTdM5wU4UQ3cnRksL+UUc3crfxI+OVJKZt+dE8ws4ek9dBRu9hO3R/fhdPKEP0aQAz
IjBhYkmwlbRJ28/cilMxGcVHhNj/SG1yzYE1vCc//ASsvLTvD0XKnvD6ftGXgtXq0CsFSSRCSgGX
KfTCjmICHlqMLZ4DDLc+ff57Y+smvfEjbcp5UGY+UiIYtgEft76x66Pj+gfdC9tVoSA8cGkev5CT
1VqOHgSalhvmDGAz4TmDtI6FI7SF8XJk+OlN9/QHQN3PCOxqnNBp7ZmbbTYOEEA9AZEin6m44jZK
WibNcsx6P/oK9tHhs/To3Z8907kG+TG0SxyPz8gML81zpbzb7G4s+noRyOtuzuONn5ydIFT7yBO+
1SFXKrxlGYUwmASr4sWuM6ZbyJ/vZCWTEfKzC571bVog1atYi4Kd1Fam4MkXz+A+TQTBvT9Ah4Vb
xbk8TqD98NC7MfV+eDD5ew3cR5AE/4J+2G5pcLCzRMLIlE4HYcmhsNFnUywaPHbDn8WoysAjgqKS
xbtR/C7cK0rrGdnaZjbvv3g3zb9SMFRTmOzq8g2WX2jn/6oPnIpW2WaQhQ6VKiFqdMllOuOVAIG2
FDccfnZJK1MQoX3fwmnDsBqxzgf/2yW9+iqgFNWhWzlPmSRSV9aGUtqfpxOEcct4H2X9D+MiD30A
kaypHfZ6NjuC8Bs93kmqUpln9hxlE59Mhdl/H3qERv1iz4TyYMJM4RpXHIQYeny7JhV7daWEaN9X
mlUcJ2kEyDnZ64x+2iy/3w1GTm+ODchiH7BiIPh35W8P79SN0XXbNtYPjXwIvdW25Nkn1GQ4P6Nb
XKC4WBR47rFaPmIywDu1lkYVav0Gg8kbhlr9AVGY3NcPxvljOTdNLMV4k5OKUxrLHuTsXoNsoKql
pu8VAOnoWGOV8DbYKA7HRH2OK5bIEjOaJM1duwLPlE49RM6pooWC4J3/NpvJSzp9ENimoyjd5Yvk
odVUTcKpMAxZbr/2U11lBheXpTtH32c4GhIxV++In9OTY0P1lW+0OGSFUjb3UxWQc+AwhEHqXu5P
oE8BcRTJWrIZGyM3ZtiTChkeF+Qemuk7Bspkq2KBNwMxkV8hTkH6RjrDRaiTUXkjvhVVK2IVsKNS
QCqxjDfcjeThaagdLnWnQyLzAcI91Dc6vgQqg1B1InwBFitm93u1I55GV31WwIk+FMw4BA0avwy/
pXyjjtS2scsOo5aztiSEva6NNt/FP0x44bRhy561X/qLngitJ7gxVX99+ovk2GK9tKKBqjl0YbV0
HCf7kcbFbuUcrHxchDX1lAUfRe5/SJr6r4QmS/VOkpYtld0WvfEibsm3NFrHUInianXhjwbmHmKB
jZYI5iogR0mcDNId3qs+Dsjnlj037lseHBHE6qjQg3t4JnMNwim7SIwrITsCYK21cKUNYTABsozE
3ghgVQklMXAnrfU4A0rhQZ1l3epdUTlzZlh6DvrxyM2s1BdTUI5mn2NZqyZXSVQMvZJvVYUt4ZSZ
G+b0EsTUNQihi+elBeakwRGZggYyHziWVY/GAWUK6uVoO49HPukK8SEmDrqkXIqeosh+WL7LD9cu
BYipNO1VOt0LsnVHjaLvP+AdOJcwug7PePxPXYd1d00lY4cW+UKtyTK1H6Fj1Gcq/HMEBDudvWUv
g1QqSxeYMp5VboSmknfqWWr9STtqII1xvKgVdrPdKdMeAKH+VsfNIdd37qQ12aQk1OUHKaCGtPzP
tyHQn9ZsaNLxxS+eBSvlgs05VF4CUGmFfOcp0DIzfxTfxpSc1fkTZw2s9HPcjJwzNiVN/K/XMLYm
IW0JsnOVUNRuhlGnekBZTB0ksKGg8+mqwNY5oaPy9HK389950IIknVJVFvF/sN0jHl5x93ak76M/
6mK/KyU2VTcModrgJ7AelU7RHYCvntSobMwdMl8QIKddTSBYNBSBL5prM+jbf48IbmvGx66lR7a4
6w4kw+3A5hdqd7ubusQ2JZ0idwMDz8HblbFuHEo2oZjkQfO8NiMaKfh6OISUnAlaLFe9A036P8Y1
kejNeNXrhYttiXdrv2lJGZKm6vB0Qo83PLdj9JOQ020atC/pyFiF/nb0KUTtX5CmuU4ZQuF+Psw9
XCfIZ2RqRBjX49urAcUv0slrZwF73b5jmQhUx+lKYmr+cVUlxUJdW+ei14d84AkF9aOJ4uWV1Km+
bwCKv7BQp8Y3J2PHpGQMFAAjxfo4G9PlwK2QKq8MI6Oqhl1jh5yE+kwni6pE9v7qEdTzYP7cpDR8
TsI2HIZDMk9POfVdc6w9B0t3YGMlaScY2D8KGu4XYm83a7dywWbsJyBcd4pU2PKwaW+cnabRW544
INAs9eOWed4EEqhV/A5liMJw5wwzgbaqekd7OsCOFge4p0QMTsCKhJG4TyOuYYFI1HXGHWvrBmzv
SK3seFMORrDFfdMxDTPT0Sfp73q6qoT1rCruD/nQBlZhDksOF7gxwSZH1gt5nL+GS/+areasafJZ
BbuFA95ODM3zkyqLPCG4KkH3V+UqYE2aKNCOAIgMH7qBldZcIcUAz/UEdy1AV5V7L7bkb6LG3woN
f0QFiSoidgzdNPshI2QRgEhv+wjI+9dLieIvMTjMpqYeuJqFolb+mtV4Ql0lkaYBXe7jNN0YO6b7
K9S7zSEkha/Ho9FAlYGIP+7KJ2+QZJyAXrKYnb/URv06JBUQXT0aAX/AU0eU9HwrzH7WWh/S9ggG
eL9VByryddM+RWwfwOeIfr3Rbva3e8ZMUTpjm1xpmK+bjyMWbrX01fDG4MO0tCHkRuEJf2+wmYYL
LePXCrjYDBlGVBhqud1jm21+YSPjP8C8ybAHNUFWzu0X0Ns4KHSzxm2rk2wmyPQ0+tQ0ge3OqPrb
XmNSqzZrTqqaxvGoSh0c0AJZrQpiUlMQFbO0UnoCQmlW9Elgnp++fx542U7Uow8huuhhKRHLeuU1
5Q3aA4BxDjN3beCHzeF8XVX4aak+XopQB6WvHXyohSGz2+c/TnT5du1LXocecPrwLa5ddc8gBBjY
eR1sGcZ35229SUU5QdjYDDz2l5GxQm6tLlUSxQsW3GB4xHcBdUQIiFvroEq5w5A3Iftr4IMjRh7C
UAVuR1K/4dNyup2PdqFp8J5VtKCJP4n5B2qXOqVCOFRuNihFNr/knjKAEYUr0Ih3oJb9SD6QkO4E
ClcxsP11KBCwJe/gY8bh5RUKfh8PUNbV1E8cH41tKG0qGIjCH+UG1AQzJ/yEuV9SqGlppXBi6L3l
D2lXRGOisxSwhXWeYM/2DIH5j/HIIWNVO/o64rPp4p9/m/1ytZJ1HFSvcNaE2P9A9TaeAdHnHu1X
S+NkhGbBGZ+ItSuTMhJTihOvlT0r10seRo/aPm0kkNJm1brYqcj95VxfMLYyfd+ZM7lUKGyq6Wgo
3wbQ2QSeesM5kBz9N0lltL0cZwCv9jKe4Al5VMwg3tMrZGxvTsR/Uow5oO9HJWyh7WCRqNLhS7v/
71x4G9FxMOHQYJzYxkzAiiW9yk1J2OKTODVyarKNTGVDoEWqwhbK6eolG9pTsn9E0j5JWp4dhJgk
OMd6PM6gqGX+g6z9SLuRILCUV1/5A1RLNXch2Cn/giEqlOSX6KncsWRetYiexbGQ9Owk15RuX1Rz
Z+r+Vt+ExVQj4vOkb6iSRuXGvjYNrT2i9Ao5H9sZF2YGkGGbucox8gZvX4caIntS+gUMXLwcC2g8
iS0pXquoMFPFrDofzqilm/APomAtDMkSNZ6ogJcSv3mg0jC8sPLVQY/UlFW2wXZGQ2p8s3sjSkrM
35RkLCLK4CjH1TBpiF3jtc/glaDNuaCppOE8egqfjDKee/rE6OIyn78WwD3fhVxV/zxaEWvI5Yij
UmwjdZ7YJetcKvlkf9MLsoTvIbzm+PRbwmJpI+9o2+J0cwCfjMgJtP6JSDs9W62MLNU2FfD8vWKt
HkYLDZDRfAo8BRwY5PZR9mxbv9pVFnoV2KVTJ8cpZ8ANIHAve+AzQyBx/gDtFrFHCI/evA6XD1ix
kzQ2ljNKPO46MAWIRA//hucpPN3cKrmUUAzW6jxm8cPTnTQdi0XM/bMGsFDdPZQ3PUTpRHNcOlqb
O6BAcsngIradlOxP52SwOw/a1aMmYUm0JdpQ/owUEXOXXhurWan59RwR55dzXyUabq2xDvQARiO3
F06o+rcnqTDT7XZ4sNXxFTaCvpBdgscJmXz3029t0imgPNeXze/YeXkeAPajQOBF0KDmGg1mD2E1
JeJWWsUn24gUCvzeAEKO8ev2YmRsqIPf8AGNL4UXbZ/5Pp1VAXgLl57UoroVzRwZiBl5lYuLwSdr
eleYd9gAuUxFk/hkjM8Y+ZXyLryo64V5B+LxzBzyFvLCtaHkWa9W7BBuyiBiq/3iWLWPtjyp6gdY
KtuD3lsKxJP6oNSSTzXQVN63ZKXLJfOljXWYkPOkKRpG69tPJaoHaRH95T792UNIqoikpg5Nk63d
dSz1tfYkM+k4SL/AoJ0iVCL5BI+1vPrurFCErfqRrmd/ezXswHfTdnlzCqk6ZoNOEJIUEOyIQcGg
WtTSAD2MOlgAX/KAbTun5RsjaZPNozEv58UfE9NFdeZ0VP/vmlbxiQwdsylsCLYKtI8Ilzm+Sp83
j9DoiHbD7XDgu07B5VbK8q5bwNdzNktDjR0ejOIVqTp9kPhbslGBzvqYng8cR1pHVOmmpTMDYqho
mS7lnEO9QhyGnNJxZG7ABd0DSwqsKwq1XPrsIH27YPNpTG61aLzHp8A5LzrMUbeORjtUWz/QXhlt
2cTrvSlqJC64HrZUCW16uPN8LxWe5OdeBN7VJAmXnpYUVz7mYu5jqQA7RpLebw2Eg8kfJ1NSTus1
eFX+24V6rtH2/Npaipo7+H8V4fy1BJvtCVazfCv1lQkGRuSZIc55/SL2IBeaKLy9EzMfM3HrU0oo
ZQczCBSNuNMPNGkg7kKftSQfbfw+I0QOEYwYAMB7veHI+S5BH9mDbV4ee9K+pKsjsb0FIstwttHX
GR1JHKWgmak1duCO3Ez9XkkZUPJNbUP6fdVmEK1z+wH1g2BjXmwViDhTb3ISw4w1UBJDQuyg23ad
HU7mFOhAJ8QHPGpzQJjaEq44aAx+m0FpFBbN0xcRqWz8orU2qd8eEsZg/eX6rxOu4M6ujmi2aCvY
s4zCD1szgVkdavOEXzuhMZMQnI0a3YZX7J1lnrbTAVemlhfwvF8R25iaJYbcSrVuZXiZBhYeAYkU
yjkz9NTGtL2W1N69+zpTsvjhKzB9vep9EMaRYNLKFQ0YntiyaMe/JUWujYWDqx2PeL8XZzRtF+0+
n52Lfw3fUGNP4dVq/OYys1h3AGPJeJ6s9OVKYRIimqGlO4R3BoBXgdRLXnH1ePWEG1R5x5XQkG4O
VdKTdopPsb8g2ec5RnOUr0jxP2TrIGB9dmIkwAuk9fYE9TZsnIGPV4Netm1DgXcHkrh6N05co0Ke
NrAGNBGgKRHTCCyKyiGEhuQQfIaHzQYYUMKtXxJQjrJe+kcmVPFUEJ2QkMqr6fUrNeUBLqlLRv1d
KwOUVmDu5eM84RYMS9RclihFeHDhanTU2yUEgRPPBp6fvEIPirn01xU3EWRKvqUEhkD5peoWsN2x
n9wc9qGHtVLb+lbeWxH6WJrw67d5I2/bZImn9K9PAhX8sTK5WP2WgRHJ647ULRaB/Rh/wOK/chKr
9Stc+HGAaM8mm0sTJD1y15VSjzvduniK8caQQtkjGC3vVI7mk6R5Kz2xCmSh45J84MzZPnK9olVy
xkiElMIUlDeEUEwrqd+jyS7wwZm3PsX4/xJduVnKEmQKYek4ygpjJrJ/HqSZhUUrZDxKdAhq3kkx
x5bPMCSayz18TDBF2Z6zN5dBhr6GrdHfKH7eS1MxYN6DsC6QEtasaTyoWdMbQRY3GhcSK2hdFVJQ
J8bVmxLiaSVLX1rchGfqfDnBZrDyodTAuROZDbA+5ANkn0zFbjIo/fYS/aKGlt6x9uotKsUgA83n
de8OO5Ziiq8SSDZy8NCfIHRFbh2bKBLVuXU7pUzYW9ZrzblvSdt6ZopVb7j9bUOLNSX+0BNNk6Vn
XsJWbUNnZRYHM0brKq7DcKzIpng9qBrKjHXSKzLhkPKadOL/dqXnaJdGs2M7vCykD/wrio80GdDi
ANPaEWWy8xaqPsvGTxAA2UXqzzq0cw+aoxCjqs4dnNna9nXCFA9o5yE5ZlR1o5VpML3zkbHJJsVe
LOVHqiC9S86xoiFh67cpXkLzZTkrXlUBLZlKIVZ2Y4Fwd2tWsN1DtNN/QJ9cJQoIp1gjJzN20BAO
JnaG4lVpIj66HeWfgpf3XWzga7/ZcSDtJhI1gh71MXDNxEIXb1E26gXqsT81fnPR/vVfkWeRrvdj
BOoqRmMQs3o2zKuaxC5VJ7dzPo2fozLjPZkjGz+veNYtD+3oRArQGmu1aPIAykXgCzk2nlPSnYux
rSXxSvAl7gOujWUdPRGX49KQ1TArGkE2zgcycuAaZY5VjGJLLDBV3HEVzBGz2kDBgLztuov4Km1h
bRQPecyfk9kn0Ku5ZqHNXS7kvCj2EjMj+vD3EVj9xh8Sj7tbw9D8x+aYXOr7W5cf7HoxZs9Zeker
Pise64zdySsQ0tQQQpB5A3BDCQh70UWplF5WmTZa7Cb1vZKXjorxoWw9GleF5xzcDzKukRU3zbrI
9jQsqXo4LrSpdC82UCkKi58TPiaMzUYtdfeSqh1HJmgCb0oDG196oz9iRv8pZwfDWeWZqY6Hrhnn
SaCxRnih90qpKW1p3V2uFcC/TsMgpf9SBszpQBqD5US3i0mTZFkk+q9FxoBqzDz/wutrPcP0Y4sG
knSt4jU2hlGEPnVTjJD3wE/MO9hv5ZmzDO1PqR+u7b59CPoXkHm9/YeohV5Vv+PuIDmuY3Knkjzc
28ZRt3hVEKDoPqDN86Du60i7k5F23NOCDdOB5ZKhCnYOsDQ1MNI8g/wBupHbhaRafaVbUoP2bzLo
XG8cJUueNjD5k4YFashaMXINoUTUSXWFrk+omz3bdpPen8JZ5zbU3U9692zjJAUGu4LmYWH5q71q
iIL98nDhywerFrxEAnSYfS+ZUkDLEywdoQU/Kv9406mtqzflXosd+iG5f0izjNrJu+sJyheS/Ziy
gY3zAZ5DKGIkxMQKr4DNcIMffnTi2SYh6eL6gRsp16D0+enNnjXh1nYWurTbt3yu/0IBv0poaVxc
BmfZ13gNa/pUm8uqlFpJtBKbGaaN9JVNEYlwMmA9GnFRVttGGYICCPO9jtEBIQPU61XNcpI+jF16
PzY7gzSUqAC3Flik6c/75muw3+IYRBEZQuFC3uuvuJJFqhJAJjS/Dmat80grgkF+3MxVkp6WswIj
qM/b/vNVZ6NT1wCXpRJjqVgC4QOkD7aLZUMCVmbL3e1O8Keh0gG0qvv+KLkwR2apPMsZw/9PkH6g
ZgBvOvypR8NOq/hF5hwnrQPeJWDAoRnZvw4LQSYPfVJ/TWoV0q4Rasmbg5vBiLiZbUH+y7rD0CZx
3kn1l0GkDNIw2SBVeqEt5zoCmriFCbkjhKB+gTcwboA55p6fC7emc94G6pwcqSYke9d14HOmL/IY
A0V2Z9K0/Y17VYCfE3xyWDVMiFMwAXNLdb0XSLhsbr6AzTPkWiF9im1gPpYVm3pLK6JND1lA8jxL
8468PqI3yjLZ7JZJbjODu3V1osnUj64EeXFaVW+EuwnzuWQIXnPNnlE3O3NlwFx7WFSD6hPIzEkr
SO2I/b1j51qPeU2iKSmLfww8uiXhGyL79YvkhMLUfGKysEwWAMK9ieyAt5Cx/ThYIjEgte6EJGee
SpmXsdL9tBteksu4ww6nP2Gku70T9rGamFanOxw0fgZfaJRYO+tj+5PU+EJfIeobcoGaj0vjQuID
rxNiXc8vVMUGUwlTkfHxhYOsZpjbaaAijL3PRSpWUqLmQAEcTXQNSXQOQjBtCxjKylF/gfDwB/4/
Kai61Vn/t48burCp0LddIEzuwZex2+49/Rdm6hyetizYZ3UdXUDBRQuKmSF3ij/GoUT2WGcV5PkG
8iqb+gsL5Szf0jE/lGXxUvnTSqPLAwEAySOo/up0oEoKptsH1bOmqPuhzqcPicoVquc+pCqVxsXZ
6DxLTceQzFkRGrepfO2b2eZDqlfT3VKMPqeo/OR5pH1sc9p6AckqphwQ9zf5V/rQ3rWFguYB6aFY
4jH7oM+GVYfyxqw4nmJ7kge4SCkHD8x4Q+vGiu6oTm06sGJ6/dXw9P32UQOl8RMcWQ83hIKvoJBk
jJDeajgblg1Tqof7aKaJ5lxC1ZHQc1aeYHmi2xBY9esTEC6gBJ/n+HER+uB0wTcAgT2f5B/JGG8L
iVEJM2Q8XgsJ4w5ACEmTpjjvjVzjGPnSOXZNvqgSxDgmUtvG0UpzEXqBQdnaRMvhW/aonZhH+VdZ
XqazN5WwLRp75iRtuw75VFn9mByxtZ09ds+Q+ciRcfaYdUgjqz2MsKdyKorGBq3nFmuhyWI0UBw6
M9VQJBWXQi0sqkMz2YuYzzwz9EGQ7HyhvUqy4YazTLDNWzBqscYOyLL8zasjVteN9LMCEUvthHUK
C6kdRMP841g0mucxKjOGPMby21mt3FQCwP1WR26wR0pVuwQQS+ZYt1Jmr+w/ZCHxzdt5thRaJwnt
GEL2myYzBOt6IK/poKv/FZ76xqc400lYYPYnmVt0xkODNepNMvNgLG866+vaAq1CDxWLhkZVHIrb
HT+TBndMltF7iofWlP4ioDlsyvww7xszx9FbfMkYTEemh4arMW5UHUQEf9SM36iTQUSRGw/+kIl9
8/qaa2AdTJHI8yMu60EC+PTRjERZMLY87pm9VfYvBg/EII8KM2Gam4DiGsXSmpVAlh5seNW6ER9k
AgYvX7DyoVXNU7BQVhlQzEOER8Ddw6Zd/pkjstfc4GA1NqHuLHSEKigPCEjYeT/8iN4Hd1eFy9Tb
nyZJOp3AQXt1QkXOC38yo2Y9PxBlTXjnTcPjyasQWMf/RufbkONDzU9/17df+DnMzObjbqfIX8nj
NNjrs555+h42V+y/qbR7aBK5xGd3lE5VxPDT1E3L0BJf1meViSmkMC1UNV6OsEdHs0HUNvtqBQEs
EvXz/Yok8Y1EFe1wS6Z1YerCZbh2lcKQ+pJGgxrDdsyv3PH6811bm1sgfHckcQwk5JtID9Odfnyj
ZfXlUrjqaOvvAKtAlaaiLzPE4dUxw9+7RI/mbWqdbkP3NiuKzWFTvtPWg7npgwbG/EWrmvGqQpKE
Ajf8BAp32RHvbZOMZxb16RRopsDJuoTLWzl3+g8naNx+Adv7jmZXNweVT/wvMKTqeW+07owfqaan
weHKQgpZJ97DyYW1N9RWV98BRVeB+Shdr9okKzC92TMRvXeIdr+okI3F6GBOnyL1BQlUhercF6Lb
TdorEkF8Gl+JUXLxmzP7NoVTKqUPchA1O6ekvDgOovKHVjRH5Z18w27CO/WeO/EdXMzme8Ki3CPs
Rzyo3Cqp0JD9yFYTr2r4/fOvINSZnsEjCxyO7/jV4GaC+fAO2yUwTjjnHqUyZZ7u57Im/6gTwet3
K8y9jZk4ZYEAkI99TS00O6+gu9rFipy6UGOrDHqsUmKUicccOJVGFlg359e74ZDGUtfHLaibHWW0
5LPXG8hLaSxeIoQNbaN+08z5WEl9Dhb/SvKTKfCyzqfECmxmrg4gHRIUhZ+KCz1dHztUmW3ffuq0
0f/66Anku6EDVi/MNK9L1LSFUjwI/0laCmR64EcVS6ePdgq8FI15GlOBlY75B18XKBsfJPEaKsJa
qN3tnafYl3mkob3zgk7uM5NIeGMEzXmRfueyXLSP1rme9fHPZ4KYCXy/Bt3d8LEd5M1oCfqAMW/f
irys+lCeduC4J6Imj2fRFSVmqXmAlqxDM97vaIalPsr22muC7NDA49ub48NNPv3t+UK47x99ZB1D
rPfHtckJRQgu/485bHLSCcwuG6Hfm3vRvl1oiwaoTcir0jenGhwVihEX35prImTkTFXb6kH0nt1X
e73WAhEI4SlauEofSbHPUEf/ewcY60gIeDJZ8RfKEcHcETaKcxJC9YogsMEbVyPPqvcuOx4JM7E7
M5hzn676A8N8WcBbHN0qlsiyO2Lhyeu053XAxmKrCROpS6awK2b8TGwBpS+V8Z0F3V4JrXpQ5khz
3kLYPEAcQvlFmUSHWaDfWQMvSCY/p5gI1MKzgrlvH8fT0H4gxVgSANklHuc1IPKf6IuYGTO2DGpn
rnDfAts8Sg12Sr1jxIWG38WFYjfEJpA4PpD3Ub1VBAAU34GUDapvjH3P0/3u+vdbE5jBX6bjMcdU
vt4gnBtp1dg7KfXhzsbFkPimDaO/gSLCecoXSCCQskljGMpEfhLo4zy5YGmTsmTnZtt9l2SJFVYO
LLZna0f9ZNnRVRZYyfMvzg4El9D/zQt5dpuMK+nM7tWwyxJvmxD6ieuOzacwf7gjPQubSknywY0V
zsNx9tXPGXiaEsqA67bW/gVGHxM0ecQ9O22VyxF0f8CO+X5WOxrFNYEl50ei5PhOL0UNSzqgf+N3
NtRaCOtr/G2y+i7i7gIXDoZbSEO8ib6D5yQ/pfPsBniT8WdhgsYocv0U0EHW+9BjxvAYEvfJG/gE
uUj7FVXCzw+cPgbFqlWMRgN4MQkvBLcyfBrKUp7E+5RMiDx2XMhRXXMoT2Z8V5llf0/pmpIQKRb/
sI07bn7Q8dy6+Q9FoKOet7iySy1oG6iZuzPRW0+Fg7ApN/UyTSxnpB/CX39f0p65rcvtplpqtxvO
8Y0vXi7HvDgkVrYaMnZ7jg36Jq5rdDVfSiwZxwSONWE9rM6wuXAHZcu0Jtg9L8ECT186LAibkox8
EBpKCMpOrGF2UqFGg7CjLSitv6W/DPlDxnZQhtUcNiHrjO3Gt77JCRPWJpL7CEH5MTSkIiVgPEJa
A04/7XQSmMCwel7DonPh/BTy+MPGDzN9XMrxcM2FRvF37aXFTYw70IcozT3NR4a8pjiqP5ZK69dw
7AjGGclrhwwqpm59jBfqHbh8I2mVkY3GBydSYgKmX1yn/mDuCf1ki4l+YQp6BrVRJI3id06hthHj
hu0tDThK214nL3qtFzR11C7mtukkZOv/doabdBzhZwzBuppF0D3NVm4/XIbfh4qKO1YpjRhkxfv+
A0WVxoavLbWgVMQWpMNKU67w+FYE7MDTB04TBQ2LZK7/71e1vBrsONx5kIfCfGmV1XUcAJOvyVw8
Y4DWq8nN2NSl9eCWwB6gXc1A2OgAth4MLaKtmwZNqX/bZF0oeW/zT1K1wxkdgbursznZ7xo1BKAP
hnK+UJXtBvKZvdO5ddmBPfZUTb8iGByhrQvVUC9ZngJ7jMpIW0rEVPutALUKk9eXXVufdSrtl2H9
pHs4IxE5aZBd0OVfsTua5KbMbSmpWulc/scDBlTvTx1a7/FbfKnCydh+E50pZiVHOsabF7Cm+L2N
ed80zWsLAiS19K74fkPnJrYYR+dyMWWbrc62peUlkQlECICzItrtb3BZj+a5GyGJgqi/nNfd0Rf/
rac3W3WWjg18CmPkSV90HsVtpmK+x9zcE7TzXUQxSKEl5UlfWigZgOTjcYBG4EW+h54q5WsqU+eO
egX54F0Gf9v6im6Dt6Z3ABfGMuDlwUebJmvY3kwr6zdC5IDtdqDqou8CLh3G8dlPdo3GiyaQDQMG
435VuLDdW+DWTbweINK2g2lqB4y0d7HByR4SD4e0zxj6Muqi6d5FleGDPrCA5xirB2EX/4w/VOeu
5UEwAhHBuJGqcJ38zFTPjRC5ruhkuH5csKZroIId3xEyi9iwNtkqb10U3I2cWD82H00hhTjyesYm
QQTNsJECWX1r3xdfGQ53TQPIlveR0akqnzXVht01AiuYdZV755LIVGo50FSmre3sS4i4d1HVYBGL
84gw5ro1HnDRwFPQ3Yyqz/M7aXE0eQEZe/1+fH7rbCZxca/rU0lWw/Lcj1KVpZXLx2h3b/Teo9PR
FZPnCvM4EnZI3LanwzrKhNWMqlOxF8ddYTj/FE0jXuUqLWyu00guRw4J3YUOOpYkK/zRfZvw+XLo
WZ55U3LQHlOR62ZlUNN5lhUEmOKpG8AaSM7Sgyev5mH2GLUKsL3qFsh9xw02+E98IOTvi0Y6z4Pb
8DOt03wY1Qz4iUCQwyB+pLiM3UzlgWoxvv7Hjow6dPhWpV3UGajv4rKdsz6RAvsPn1Cjf0T6Njr0
WbxvSi6vB7dTJ6UZJuQNzHI8BRlzwXm7zKwQ3baI7jjwRpAzYIKDOW8Tv9AP5FLlICcGJAXHPMhb
Wgdv8//J4NdjvXrqNhMOQSRoBekLPvSiszPqGRUadUrapzbFQTbz5Nb7Pju4Qp0Mj4Yh2reXwfbS
tXq8yhK+9gkPyIYR5rVgs9Nzhn1+FwuJibKXW/n+3lHggH5xutPqqlE6BpkbtdSDGrifyKUpD61r
AO5N31qR5Gmgy7HNCMQA6AgS3YidfGn1Ps3a41KvO7FV5ABcNOnOjPhq9a4m2DLqgDg1lR2yY0P/
8GA4XHkl7Am3GoroM55Di0ni4/ZxdBwj9gBLVvOdCmHaYqeQbdYQuu3PsthVXC7Ydb1cUYKobk3G
/8ebJT7dkZhRhoEyb/VQgSJqJ+W1lQ2pwFf4xPwxQdl34tVop+1jDuAVgfoLiGSYuHDGKOQH9hQI
egblCrXCn95PqMDjzhS9f5JjrIe4qCG6Vb+Lyn3ZX+GLns4ZkTdEMPf1lxp0hsI7vJUxR+fQE9m8
To703APAZ8vLigG6RLFCcSjIsqTzvTsgT1NvWaYoZeZtn9SI1mo/9RrihqfLvXzhgMqmljlEEPgx
lsyljNfw4XCGKjjGkYXo4vWIsAEHh7tJejh4lxIiAYluKn7tkmZO50PGLdLVskhpPsiXmZoI4FRi
qawgDm4pjC85fMEsgRoHFfRSwQnO+CH2iFMPJk/079XPaEbdqTxvenFSoxNquHIkO1sD4qmX/yCs
blCzRu4LWevYYshdV8Ccc5dxuZ2rKxhEw5pQhjKGx0qx5e7OGVDp6Z0IMKOQ28KgPAnTQVOaFtJm
6oLlfE3sOvNmHnNzUDrmy55IZ2zU+SYiPy3nJwPgMnHHr6im7ClD5W0+6IKjWKPN+xHD5RD0aypE
zrnjGNXHBdYHm3hDFnee9/Jv/HLgV64m+m6B1FaGSrfHYWtdsizaIlAx5gf0sFdUaKGVNBBK5pdf
xFkPQXxJ/hZNRpEe111Pw3OBF1/4c6lKNRJG+FifbrsXvgpt5IbeVHKGw31JeOJc70krs5ffezR+
t4yaEQWZxgnm2aRNrVuTQNGG0oM36lsCXC52JaXBvkJIqv98fXrfhMyooiKjiz8/Q+dfncJh3PQ7
moid9GmNrDGylBKrKEPxBWPjeIGtiMJ2x28fHPQnlWnGGa5+EwO1fjsaU74OieMc3H3x6CYFLFZE
eXAyu+eF9T/gEt/WKr+3SnlcFn2G9inqe03IHWWqlLZohsbI6Uo0IqdiNX6hMJDNpOXKZ6Lk3x2c
CHwW05blNlJ3LfN3m1K5BbYBmkcDTdjr4T7kweiOvlO8SECzipvM4RsTaR0KIvd40vQJnem2epDV
LOF9/NKxi9zl9H9cKtRRphhbQc2eAzbEl9ksTLoSiUHWWJ1+3O14Y/yntaSpq0q0vuXka1krbVTH
oSuD6IWdGMNxqTIkN+ga8NBMEIjha4+/qM/mlSaj6brDpYTpWfHEsrfIid/f5xt+uUyCHBGv2E+b
XrCur8Ju4WrH1TSx/DV1QLj6uSwPo5vjtk8KeVBCTWWCusHn5Z0zl8+VYLfbuVTJ/sBM6nWjHpaw
p43ZHPKXmornJMV4MbByn+26PgS9gH2wzNiZHHm+ufBLBIW7MwrVq0Jo9Wh7uLYkEnIhXtqdebo7
RMyJLn0wSQleHqSOu95XaLyVzHORZAHavmpTOt9o7Fs1Ns/igPUGJhoBGrASTl9zsqjHKr/rpGMt
zXLdB4oZupC3QATMb1QRl+mCPPS790qqr3rN04pxgkLW5ASDfCK2NlrJ19FJD/h16/Xt8TQk8wkf
wqM+USj0wDuktbZdMpm5vpAPaocnBD95S+hnxcKFbFuLG/4g/nk2E7PU2b/IlMkJdzhUP56n7c3Q
phDOvmDCZYagwbYCGFeJt+jgVSQCFUNT86i1Zv9sUseKdVRv0Y5KmnrpWIxq8uilAQCHZIakLaWg
P/QCAqoZUT+zirDqbFlTMGmrg51FRX4DCfqjdMpaDGMoqYxV4iVaNkHGRMaj14bJaE1EJ1pbSTp/
8skmmeMCqWMlFEk6RXcFaErmwRU4K9J/m00SRahC1+kbYrp+G4DR+n08siF56+iSSdwmZ2frleix
wdpjkKWhPwaRlewQZcw3vw1QygNi8LCMpRtUR5bz1obWmLcDr35DOWXSJEp0TZV6pyieK/8p+SiD
8evATkvLQufxDFRCulL/gJljnxmjthshrDOrf4hA9k3u7bH0lzVOw7LklclOODfXG0VnvbuYQJVX
SX5guRZOhU6OZ9hgaNRHU/dSyny1D7YdtMWIHp3Igi4Jzk+aq/sjJb9sLwpq2ScSMwWQr0LQCaRq
78cN/RS1yy3paScoAaXPhhHD+9Gf1kZnyQRptor7gqdEzX1VyZQC6JrxMo6FIhklv5/8z0imuKEL
noVUKQKd7XKtb6Rd8gb8lr5xcuygjQJLP9Z2TT6hH/ve49eCEJ8ZI2X5zyzYKUiD0bAla3CgV7mC
WFI/N5f9CVi1I8rdynORWybIsJURX9o4uQ0bzI6p8WwIiud2dJrYc3W8UyG7fneW98k0R1TyyenF
Atk+RQYoETfSrT1VvY5rMCWdpY2GuCBM5ybsYE/9+WUVv1sLCz91At2WXbjfFjr/8zjBMTtL4aTa
zSqMEBQssr/oPj50GNc8eytGQqqqo0QJjj/Cu1VSRYnGqI3ILQcu31ZyQRI/opXu0XlZB/Xm4Wog
7Ua9q135AGOZhRK7rZ3PrqNsCstd6K9xdmQwJZ2NHvH9gkqkdrfamviXWIyykAwPOm/omqS4n+fF
xOSgBzYUEjX2VQXOiVNrEw+bBGwv2a5icEas30ZJUTX3qxe7JVJUiTtYdCbKSJQ6QAz+m4Ls2MpG
zGhFnEf/L/kooiwZqC5DclVK0zGIrWt+6Ub1nttgAChP/6HZAyb+599I153jL15YDR9EC/By7toM
8VVKoOmqq9vJ2WIRFgJyiX08Gsau2CGEMg2foZN922AI0Qc8A+74iNlG44dS1b6+vJQrZfslO6k7
pN3PnWm5fFY5LD0zx8MKf3jUWeMKRApIyllrV4OChfynNVvfv2ozKrWVX0+tOYbxWLLVzUPQdPDo
Ab3iK3E+r0S0ARq1Xqllkp1BW5lOqBwBbyZw074u2ogTTZ25YxuwEEXra53rYpg/bkKZbVpILhbp
c/FR0dqdey9Rr+imHGB+QJzRwPCuNiey5qAdz2bAFGl4aCd4lfJyf1nLpCeV5XeN9hfo+mdO5UTP
0xmzP6R9QNHk+OP9S2MGyV5+Pk0QO2FLEEpgKfwtDjbQYjuLry4BLzjefd8Xa838PPua9/K3gCv4
J51vCF7JCYM2O/qFtWnw2JUh26MlVEedSqXxf4TORs4Zs436LLUM+SignO1QBPzIWPZiEmqTem0q
XAiL4CHqXSymnElEvhTGaTKwOvxNT+c2YsCFDvMzODVrwMQ9/ZBSB3TbqWvKYRc8H1Hums9WpZSf
Nf9SKJTNvg2j4bNZpA/vtLs4zeRIdajyG7Qh8W83ecYww67BzihgpvsXusL1jXX4GMSmPhr5wshW
D576EOH7PpBPLqKTqzXWCtiJylrerlAucd++0/Yg4NJyJg1BATVb9Pzrv/YDQ27KRuDZ1CgPuY53
AoZnzWI2d0dncjwoGm+X/y437SX1lOF99+xK/+1X9G6xKFokDOJCH0LuLcpKjRWMMNZZ5V+k6PdP
GtLEAkZJyOHTqjUHsbjqf+yr4js03eXxYYJtgku38LZosWoa9fZl5fJUFDef42kUCFqtuwBIvcDF
WsJsJuMU9M7wXB1sB0OEjizXQdZ7aMod6nOjefJ3tpLFwG9p42kBLXHn0IbiXFxd4ankrPjHzstW
UMEVLiNS4sIKo4sTSYb6wPIQJeD2rPTXA903DhVtGdiLsF3JmuydSPpvMTOT1qm027zuQKsMCupJ
SEmig5H3Iv2he4q+vP0TiMkZukKEPUsD1zL0McQWc6f1LUUYzuJk24ALO0UUddnZkRaF4Ey+3jtP
LiNJnuGpP1w7QkXpg+VEV8jbOoFzyIBTpHOMz6tPkWkkplvqF5sEacVR5XyV9DwTIjxVrpaCuGwq
+fQW+5T4QkgPIB43qCAJW2ZlkzdVfZdXH63T1OjxQs9H05sVxI/WC/nmSoOVVBOLCH/1OZs4Ul5U
3thWGTLLff0zhYA+tnMcxS8WfnGJM2lBAJRrU5jXURqel0lLR+NYHz6tQfPrfYdsIsIG+N/KNMu/
27DtixO05Fzdv5QSIgz8mLc1rMWxXb1QsP/iXzFboe1Y6XfrRth1fRwcjfM/+afsb3jFMJ40g4yM
cTKzOgqgPiDKv8NHQ8pIMwkSfXjWolASQZd9yL4oNsWDiKG/vCR9ER1OxCeYeEQQX6mpnG1bH5/S
ZgLAqbWPhbiSrpsa/E+TfxEULZJ31ampu5sefScdbLZ0tRaLJK0NbsyCXe7S1rsaMCGYGhtqeH0S
5VK+v1zSmz8ScbexPx4hCMotXoBXXs1x6W72aVHoBHyOmm54xtXzinhSwAx94ePC0zybIT6ykBWg
FxT3AW231VhSUgtTa+UwzQ668lQJldEtV4w/dromz/KsK89XkA0NwValW/xxFZtb9lutca763nvR
vavsBFnqpfXFsbYr4hS7yCmhh4LRTd00Xu5jVty4/kNV0mv3gUX5RXpMElcMxk4rm6w8O7g8YRT2
WLPCg3Tvf4RBuRQeaH9Ku7YEA80wMnPC24O7m3l37D3tS6FH0As8SeGG/Xz6lilJkT6wASanJT50
V4gt/JQpK6O0TDUSamhESvoj9vw9FKnyDITtskUyDtF7FGy2494ElNMu7V7XFfM+lANEyAS418o8
x9Mi4dFFqA8/khrHYJ9BuoDnMB51qRXRc21oU+wCFyT8QHoKu/T03Tnchu+xKrjZVV61Eh6VOGNJ
XtNxXgJ62hIo02H/OMmNldo6oSUvbHfQra4om7MNMo9WgMy4KsuCUoVJPkH3QtIdrVjqPLQqqktZ
BSoDZZ0hHfj8TZrSFanSzZahrs7caAPoIDTC0q655kvr9+gPiuKXd1iBttTnMHt5lBixlHpErfe0
aai2eyYqFobp9sZxAn+2+4UvZq4MkBTu/7ZIa50/x3LoBOUxRpB4KTumcmhNuvXgvQmtVHIJUuVX
cURtYCdEMQJV8YmABT6oaqV4PRQOqaYVXsIVEoZkivteFBeFfY/cYbQ9p6L6v3BRi1XiKoz7Leep
Zf8Nd1sEy40mNgSib+qA6sngeGJBQSR20O9ZfDZELzYu4yuc60cbx9VGE3wdN0QtccXEriJNIHUb
03SACY5PM5RosaLEjcpp2PLFwsdv48WoZPeOWGRhzM0mj08DYM5zJDGg/26I/QIpqQaUs7YuitQe
9C8NQuPiT7Rlk5NMEyM2JiZjmtxdxWyRuxLZb2w8Os2RnYqva9omczUcnPfYaJAkHD9ewWKeDn6Z
J7yPhUt/3NT/NGyH5tN9Z+IiXCsI3JF0Dc14youyP577g2Z++a6XMp1zggqRIVa3zouc8jIAAohR
7kZjvNyF8BgtQegQ1fNGX4S+uO2LLkjGK4jtXZiOvnHjuN5AhXbK9EfN88aDc90zcziqYsmUuow5
3qfOi/bWm42G7aRwpHRKjl3RAlzC3rmaLjs54L2pIva4xQaa7mkjPvvVOjgfT2DQv8SP6ACzDe3h
M2lc56slHxCVH5IWPjRP5FWUj0GLeZ7aaRjy6yxKNJ1aUUpkbnicbLDak5hduEJ2jgkgP55RRzVZ
CgvSNcfdO/JixSiV/CcPsRfYO3JSudd+Tms/RYCWT/ycbBCzXE7aq8agI24KsH/w8FbKIK9/ifTn
Gbp2Lyy4nbL27eRny6OlfKNtdwWkzEWDghPjvAwlncj8sOLULhm7Th7s8AdyB5exE6QVaZ01CJFN
K+5Zi8HBOcqJQfnagvg8P4wiqRpcovGKO+srm+QQwOcrTPlEQcYnO7qsft3y9O3j/2lacMM7vRdV
A8u2Og2OwucMC0CgChycXcBJPlrrFF28apqBDUeOThhvfEegrTNe2g1ql5sT0FY59FWunGWPmk3w
zfEcrX1K3pgkeMS+cKbKD7cT7bLv0i3s4vK6eW/9gCM2VP8Wg6ogJ2c8j56yD3ujjeokkRrL37Ma
QA6zy/p9khvWbfa2If+hHIyDwkDaCZEGrceDbp5x4xjvMMI1uex0N7nJrMROAXfaqE3rGDhkhjfZ
nNpXDSHGfkqTAbtXCisc6g4jxMI+IJJxQHaqi/0wEqETqAb3l/Prmlqygx/eXN8JRYoC2oPIXJHD
T977vea6MImr+UVMO1+IYPtYo7LmCXuZ+GL6kCT3B4xSMN1jWF2JdZy/st39pFefKjyMzXg/6dl/
AAA3PNJ0IeHDhNpCGn6hFXMpH1xDPrBPgtWEGLFx86GDwtgCdAszq0s2WsK+aqla6jYz2L7S7sTE
ftD+IFt9z4RvVKt3akFW68GXnQguRtGVxt+IjDUyARTR5Lhrqk5pzDznVDUrP1RYZvmpNuEtvN1B
KqGrE2Qan3l4sxLZRju92W5quXTBXVk6gDZ1e+DXoP9zKRZouYQWX5EXY5nSs2782eIbZj/wBBaT
ILG0hmFbQPCY4y7M0f3ftuz9bQZxnV4ZEVHMuUJF3dwlQMCKZ7XTxsI2CTdZjDZ55lnX/VitdxVV
HlRe+cAmZKr7IZYs8gM4Sx70ODBvpZtEcm/hbgOtWCB9yNeBkBnSyRbEN0OWzwKjn1ALEPVF5HCG
NpPaPs8qepuQB4wzMXYxOH+w/Pl2iAtke8/vg0nKX1BvneoqierJa8Y4dJtRF4j+M+Ecxt47RHCv
xYoe/dFDjr68n+NIRaYaaD+5WuQqjrSSiIQMevOjOEqwf/02a95udCG/coWKO7+HKYDBuz+t0ChW
HV1CVqLwZjJdsugUQfYCQnW8jnnMuiu6eOUnJNVf2B9aMoTRv86hRyMOKohi3YBF2UaGKTJ09fce
Ol25J8IjGv8RN288O/CwLBhbYUo1h9wVn2q26GiQYYEc1jtu1gtoDtlDAJYYSLA22qTb+3zMF41A
DAUqRKiIr6Uo/6/5/YR9kq578Wj51KiLseFTlQZTv6nIWJfuV7Sw4w73TbQrwvlKSfdsvJLvBXxl
UNgcrxbIMrm0TkkHmjrtgdILYzv70M/fODYh4avrOMiiuVdHNeV4VGOcAjYFywVJgAvNycD42qGG
Kvk4ZwU6XO4mCPtiOosfC0JMfZSpTkTzVqG5qgi2USlrAiRa1ICqisPA14hfGJ2bjvdM+RjWs+J0
JzgyKRrDjnpe9yEMIDsDjp0Sc45cm+LDDK7zI8u+lJRAX/bz0ZwMS6hFYOGP9ZDKx/KuLHn6VJ1n
P+as+13hqmDKVr4EhJjMT1gKzTgOwLtnSlCC3of+Q9fJjfr/3Ca+Fp3b09s9/nQZ05sEugYU/MUL
7Q/55tJJtLbWsVUNbJxxCDggYgKXo+pPGhnviSkZmHCegPcOwiiGk0RP0EuG3W1oT0p7B5GeezdA
JqqtXVSZI2hj7F6EJwScmDgQAecJQ0jmhYfQYkow4wRAu0c6BRYTwoQb6CC9DneNRhAMxdDLhcSX
rIvQodEAr80H4GkA0ew9UCuRXGD5qFGsg8BX+AhIUjiQrRK48fc3WtWiDYRIa/hhh7VrSelytIQm
3vcdop+IhD02/XB7tQGtMhpqQ06oHUOCT9jyxdQ5QRbyd+5tpPRWXnIMzV3WAQS0tPUYuF3nGGbG
Rsm5nj7DPsgQDYMskZNMeDmnaVbRLbXWnylXR0ruOxZ4I/MLl99SQnj6EdLsZwyNA7WFFN6wDh3h
2XaZRQ2lrC4JDScgH59YIJEU6RzKsLfsl5UX4iC6Usmyj38T5/b5yLRSowzojp5YG4tt1K0IHEyN
hKAMBUaa2IORrEIlUn18rNItv/ad+v115kGHym7mt2189+1lDmFGjRR/fKmSIn/C+/NIDUGQkS1Z
c7utrvOcU2di+4gdhQYj4I0SSaLpqQp6tx1Uq8vEIGsYRGzCDlYbQaQ8qWArpSQpl46qfWX9DN4z
TggZheB5AKRmGTYAOdaZWYYvaZrQlwejTYAMIXa9Ch9VssG8/kU0eVuKs5iOAd5Cy7l6xhcRh3dD
/5g0C5UDQbZvakb72FFyDP9jDnvOd7HLKqv+/PYYAOcEZwm6ySeo/5jdTFHOjAog7iP3H8s/b3M0
QDHIraGK0E27kNM7X8rQBvVqgyPW6rvy4vF/RXfbiWL8HSTrUnq8t3dLp+3JMvQpqDM6n5nPLKW6
TQS6Sl/Yc37M+zmLtRgD7S31vbiVCx9DQWe0H7PSpO5pAsi4GkQmSAy2nl0wLjhMNQjd8wF9Tx0G
IPSo5NpQaNhCQFn3krpl7beyKBxM3/Oh6stZzHLwZntR7VThpSqrPvnv9jpot/1yJnZEAF2wtgbE
qXTbnErJxldX2W+nHG3hr045mf9kY4Xorr7RYQzzSo1Ocado4Ryvzxxxhr9Sn5Q/TlcFJJ/NIb9z
JAYChf8BDgbPM4dq32IhS0mRwLJtm7oijBsz2P8BrjK6cMSM7pFdcD/yvOV128EAdJE217f8mbEi
MAPH2YKEDXyVIsQBcEYvqIgqdRLdePPze/mnbMAnzAQp3gTwoOktOH56U6flt/7zG4oOli6LxYHh
9xR+ZPEpT134NleHOzMAtya/XcBR/Ahxppl41XDTj03ww4eFE+LCG3T368Vql0ZvXE+YMRBMBn7w
mvCpAJKju/qgQSM2o4druBPbkzl3kpZZldepx5yyCjYFl0Z0LXAusG221mWi59Wy8xQwQPRltgYm
50SNIR+abvLnyz+DVFEf4RXkAKss0jTmiag865arVS/3X7bGyU/inuxvh9EJHrzNlZXcWkkcrhKd
47Sre5SbhSAN/NB8iXjxaeRxM1gthJcF6Eoz7rVjbFxrDizbWLygsuCvtfgoMSo0BWXr0oXeVJzG
jTiLmW8+SyM+tZFlnIn0vodA5lsEUBfcyELGFWZl2+8YIkW5EbWiZp0JcaWJpnMiZ0uyAStSNQXo
w/xW2LWlr34YudpgsqjfqiFTDD5Dbtju2+NdeLmwN+ySN9Xq4ifJcrA+FEX4I4VAPI3YrVaVY3LU
SIBKygCsVEruK1PcE077YiaAh5C2sCly8hJOGTab4Tv8khLRtdnN8JtKl9M2vK9i0znTGaOx/O8+
BPbJJ/AUVwYdhp/y7dqbXyjWtRchX6HkSxxP3I3wb3ryZYHOpZ1MWpKzbDP6cxoCLS0d8wtEbv0Q
KrMZxJulDecaJghXnxobTmoTfLwwMoIQg7bvfuyg3eudlIVqCZqAW+EwODiEt+l4WkawNbMmfDNz
mBk7KqgpVNMuHMxH3HLN7kjhRhwQ9thFalP58OTELAcVlsZ7yBXNRcBZgjq92Pov7K3rc9gy5afA
ga+zkEZf4gwGt6W2qxJzBbTYpoB6bWR0bOsHfUEMTXMYpZzYkPhfm9r0qdFGQd1uOdSREYDmMaCT
kk6R2bfV7k/NZ2ZPbwlS51Gp2Wm5CGbtJGFgm9CZzIYiNW7balAb+ICIjL5z3etC8acvdpqTXxO5
cOZm+wS/dNftOdCIo/ixmsHbeGE6YWJekOQotZKBSXZ6s/UraOvcVJtCUw1npwERKliCluEa2kez
3TfjJLDdBlrHfgjMyQDmtAm40A0ny1cQVkEJ01eP+fiazKyJMDz6li8r4hG2a/hOEPiMnP0M9ASq
1PtqW+bjE6N17vYul11zhdq+6k3q9Mz2dWHCnyWrWtOhHQq/8WDi9gpK3sSOEitj38p3cfdSpp0d
GSMMnWIyTIe09TRtDl5b4bWRL8Efw5sTkIhGh4B0xVNi+5t4jtXlOYJeqcr/tT6oL2T0FYiIZ8GV
7Z4xVSIQxsmKW60SwylncMkrB+RoEYeBf3On71alTkpcwY1EksWabrigOg6bZB2gyzt3PaaGkKiY
37ri3Ezz1AVz0kc0E1PJPy4SgUIUA6v3XcWBSI7eK1dBB6fRl9U5JtwerPn77jXZaznd0At3iZbS
P3SYi2Zkcxl4ivBbzv2bMjYUi5hl3XpCgmZiuwoUuo48kH7unli/a5feCqoZtn8uMm3TM0S6ShZv
OHoIiQ3LzNn2C7InQM0hWtQBIepVZCBaXm6NPzyuCsD3HVCT38bpySdkI0w0U9lqctQTmJJ715cJ
z9Vn8O9ouqcuyyaAoZb16YLn+9lHJPvK50x5dypRXjG28Efe+o7kaz/au8jCHzHJYfvXYsX7pDhd
MESsdaUdUIp67/WFzmpRp3SSVKXE8vpHaXF7ofIWKKokcRQjn76MUfr8Z/eU9eFV5T6f0nfB5J1k
0U+XsptiWI5YiXI8cO2tgCt/EudBHl21FKIZM/FCMirdEZ/kZAceyTEPX864EdYWMek5Ia0apf46
5UVx4+vGNqolpBJvPkVMAsunCoTJ49tJ6G4jW+/I2MGYXdy1JzBySXFlUOvQMKNGvixa4CypN2W5
KxVN+nIknUazBwiDj35kRv06dMn9iyNCDtBTqYAXmw6eGa7FqhYaUCV7iwf0MZ/sDFQ+uz96devm
igVSgVvid/mOQFgMbdRgZ9LUR96BUVpwGl06KzlQUg7AmVmWDM5a5HK7kH32vX3Nxxjl/Jku9XAv
MPpbrenixmCE2VvuP89uEbSQSmqhV1fGKgtvTQqXwVnAONWy5GLpWATXunIyE7yYjYgdAArfKsHt
fKGKofmX73t/5XVE6AV/vvTMLvS+YHvWCTGCuPoM7Q0rvcXUQd8C2xwkUTyq/mXakLXj3rA+OpbW
Lxos/m3DYR2J9DzQoCor2jCwcU24QThueLK4/uDsZ/P22I+7NRKKPKi1b4i5yXzbpTXz+57r3zjy
suM97EZNBHEhDcHUl1+ROMCteSfCT73lXKRUETqLQnNUEAhcbWC9Dd3Cr3dIYXTOTuQm4XJOivBB
VoUVYoMlk99a06wEvIYzKoYtKJsag329u373OY1+QlbQ5p+UsoZ1xTP5t83aQ0MqaVoKWaScAX2l
R7JVtnvtBz7AuKwOWFphyMyDcts2ofcfYUHC6LcB5Yu5IXxUuVo4l6swh0Y8Kw8Mk8QP0JsH04Ng
r7g5/s6WA37rNapzPSNn9gwUlcaYU7E0Rbbc3eQ6SY7QqWCsV29E6cfc/Av/qVJUXz04Rtl3eLSf
g8VZmPz/0TZJCfkJHYjXT3z0MuOtrFw8LyOOeA4uPxmqGqf7K8TnqjxW3R1dV4M0U09OdRhF9wRC
uYKWq5YsE8nO0QxkTtS8msXWsI58kJ8Oe0NkCDfd94rej7WtQQe3yyWf4nsPe0i1UYDyhANY/pSD
phauaYohiQz5lAuIF23TgTD5wU7Yg1vJEFKyKigBxdPj4E/5EIU9S2QZ0CG6LXPGAUbK93pPUW+N
9plVrmdwZhoIpS8EdBzytPLStU5b1ikKwTioLNQTxHKYQAv58crF7RHfOzZT2kTEfMFTcQLu2+a5
q2otV0DdvWoGNi8s5SZ5aXBLro7kotswIcvf50hO71SQ8XOLRrlTPExR00mEQDn46lMvrI3wFAkp
+oBMn35+aE6hQxuV54S1Y8gzhY7hsFIX03ySyJQlgzSKusjdGXDTr59cJFg9faxTIDDT61SnG/Nx
tHA5JA1kj+TQL9vZDOYQQH3VNB2+ve7Bp0udvpqjMlPeJOiTzoyqzjXNu6dkMq+CVezlI1LRraY6
r3c0+/d8ePexqBKnNA1hQ+iPUvSZqBLtdaCMtziKBqR6OVyetFGlVeYFyLBX63MLh2FZ6K5QvSxO
Na8/ROlmlM0F15Hu/4SJzl1P9cqqU/CXiVpGTO4kj9gZ8CvmKXfC8z/kAG/tFsS1VrFwyjPDs1Ec
84VehpneJ8w9MhVXUNxJb0PRKnkL2GBkqh0OGT/zr5XeIB/SXaBwfPq9FgMK2JzSKxJihyp/k4M8
mvGpbpV47Lr/qPHMGzs1kp84DO+lYBSlL59/i0oTgEWpH+XQSpH9SnXsdkZJSg2Xp8O6m3VuCBwq
I4bkktVkNVbfOEGLlq2UwYtpn1co3JaKti94R2YkfLnXj4Lux68FcPzYOV4FTbnjv3H6Jw+26TN9
IfSd2wndV3Mv4GnGWGnN/tC039b2vm7xqejdl/uBklWMcZBpTUgJdO9kE7YfDoSjrAWb71cBUUcq
b2CgAxsAPRK9aHoGDuk9gAjVABI1ErlG0CUNcDNGMNDdAHdvgVu8k9KXB8osowXR/VWDMYbgM4Ds
F4BPv+N/WiBEofqX8/gyJAzJpOSueKcC2cjXaqWnwAMJbdHbORPALqf3L6urY50blkJZO3XqG8e0
0l1jeFTmt3P3JRiMt9hE1RcHadA+dgH5zTEXF5e9uZ470nfcdpF5pWZTRekxSvg14x7uVrzoV90v
JqFpm9317CS9hJPY2tL54LhbpgJDBMOmeGsHrFoGVyb5nKCa2R7z0D47SykQrIzxl2vpD6nzko8w
+++UKQivyffAzbZixMod3JqFElRp502FSKy2WLTqBk70MV9XYrcaohEAmDWaSEwEnNrIgEqzJtf9
PzLR2Ib77AdTTkNgBI6sJK6RJQDO07XLKMK7ETgz8+FtgsjN4D1nx0VjtHHkq+ZvNqtUlRJSb4gk
fyonzjAUuk9VETvOzeKV4k5Q7dnq+PTQvZhBUWscWW/PLoK64T9zOeK9Dw0bR3hYXAxT5DBQB7Lh
tN/Mjai5oZXCAH7I80bxTJ64WjPttowXKywTF+kZUu35+vXTIP1hcwY/YpTl+S6jMc53av10WkpK
DOVFRCZPou2SuIUn9nfiSdp0m0C6EPQHwe2auE5N+gynyG4EVBUDGNf3L8WSFGwnPrfnYLQoRjfl
tbRwM9LvcStpHmWbtG+Hta9KYRRKGK6tTv+warc2EUqDhwUtWZMLGjUscoFOmOjUVTvD+pEoHlMX
o6njO8JaPYnYXaE/2BiozsOTDnJsJAiD6qUDw0O0o5zIsFcyCPfB6bkrJeeGIzuQibicBVLJjnf9
C3C4WzWiHNBszSALc9x57A+VRfrtpdB5eF8VfkeXBkzwFKpM/x2wprgiStreBzQnj1gY3/MXlf4y
a76ZxFbU3ufIvb1YEOM0T/iqwfzMHJ/zGfYpENAyWt0brV+Yd4XUdUgQp6ClqyavAbUYh5kskmah
GpfIr5DA59KoyxQryObyWVp2N29YDqa4K84kOcE6lBLniKyv9v27SRihLO2m/eWnncJFG6ictELH
ifphNSAK7WOLpNPaXPAXNpBoBtLUbkcmV0G5u6BCXjIKr4foBzvAbf4oNr9pyFYf/KpxTT2FafXT
ioNCwsu0ag7aXy1MgJVlyHMn+5Rx7VldmYsprdssRO+xME7zAi7OQsrwrU1JXjfOkHGONwOL1uiJ
I+eUBinhHR/3IIoqcwZ5wYXwzNSjHwokpxNEqH+ZNKlCRKC3Nza41pblZs8/3sWO5Z3L0MOeq2vg
KS7IAroKZiktTZqlqOftDRgoTLkZLY8EX/GLkcDxiojlQA9yLYVW4YNS/wgRJfinR6xeUt9BUvNF
qvVR0XMvkp7wMEAm3ufYEDLJMWpXjFKoKD74NrwfKzDhEJy9yifUmZa2Vt4CgeMxWHpdo4jJtouQ
PLQjGTHclguQnMIhy6fnP6e1yGNpR/PJK/bH0Y6O5w6XVAcJa/cwPwjadE0w/XqaCvj27SrLimDs
fqOnjlHL8d75a3nB4rxNwHFvy3sPkUQ2F498dUUh1K/NzC5DlECbL4NT6WJxdhfblyd2vOqCY8uC
XDfmq2G23yz9dYCzOpUxL6u81bM2F8eZIexe67YbB52N9u30qMosrmExIQNvKMugpbZJsUxHaiBl
gbMN1M2fhPFTlio3O4ocSKqB9+2efopB9Avf83woZRtIOaRzIF0bh3wkHxITkqFsrBdUnxm6DTHZ
VRxrl2qAZO9sbhJQmIvsLhxAt4NzO2y3Ae/lZjzIx+vewImJoaMQDR93/OAhzaxB+WPsS940FUkN
/VmB9jIbdFPHnh8WsyT+Z4rZ+1Nr+PUmxp0WSdQtyHq9hZuWMbe4mak6FitqjFZHHKDostKGP8Yf
u2jNxeJPHYpZMFOSKzy2ZjU6BTCLmMmnZwXGpMaejrQ+hoElsFfEDqRohmn7Xg6eP8vSmGl9Bw00
ZRkT3ErBhBadOAwrDKTGkKLm7UADwVCZccFGW/ddIg5fcAPYKYYfATfRHWj6KZJCb3/apfUe0p5d
mvtwxT+zAgzcFwt8yDtSbeMu7ZZI3xy71eWixYv6PxaQxiXeQwphOCwOcLOPBnFKpzw3oJqAVHXi
0hECxhpiCmDWzvAvO4IZ+IFl4lSm2exvzSrpldEIwuRGWddXmP1unGzz0kYpif/mDnPxAFntC/PM
mU1jdbkWvo3Reu5MdYfBWMmAZj2BShHtACsdjEEJPKowddYhSV1OWcHh4b/W4G67jrE519ELhvnl
Hs/LUtdK3TxGExeuxjSoTSUMsxaNe/LzscbawJI57xkc2xpy3UTg3ZyY5CN5OcUyJaZumMQnczlK
a6XL3C/smAzvEd5pCDd8oZsMucsz5sRAO4UguKYbwA0nos6DVl++YL4RupkXD8m82s0ooYJA3YJy
zyx5l46uD9eqLnqRsiyvXHZWzE15RJDcaaeV4zSdK8f/oSdqxqA4cKWtTChk6JWLv2fyy6+bSLh0
oWpFjXPfcX9v/OLkkf20nYq491qwTovemvIyUivjHoNN4hQ/V1cS1Mgeowi657zIkDKNBuQWC/6j
PNVa++gXhnks1z0oefhJqd9WmwYLaWM0w/N6VSbCa260ElekP9BYli4y1xPZUZTUdmuFeHSo767O
GrVGAQXHO49tGjcORWd6+nrd0RPEmyriv5+S7CUFGOBm1wJfgCVLVoYQPMaY4SorhZxoGd6YD1pW
+s+nHMMwV4Y0H5iU647A2xv/dBpjkyVvTn3Likxii7hgOZhaHuq+kaD2OpnAZxL8Hbheq6n1IOxE
aFgz+ln/a6QJTW9ih4HvGO3Mrci8mLpzwfov9Oc0BZSaKTGxVS9maTV1+E3hZcmqco5c2xahtj+t
SNdGMvKYnAQJFhbai1RlRB0s8P/fYXjBXLjOIDxktdm7EIynL/4DVhxwK7fA+QGV1lsLfM3OQCDD
Jvlx9RdtP0As6t4BDg8TjVZKfFtDH8i4+cw06KdEP6zToaGjHNAh1bZHqXezabdCKJJd88Zui/PU
jQMs8T8wxSGkZEXLEbeZQXtmOKTg4CPmX8rcjNIk4GEUp+4VP79yTGEt5zIVeaTmpNo0jmTYfjVP
yNdn9oEPuKO1vCn3O2NWhARqhok0Mb4VauHV1pTGQCkl1nPZk294pqQTf0jla2kN4Kvd70CqC8kF
s5mWT4gUElMAgczF63e+S+FKpSzq1DnE0UUfC8RQjnMdpzLJM9SezgrJV8ix8n6N0yB66sUL4dzG
IL82uMxW5pKL32Nacyr76H+U0dvdQiptN5dxzYD4O9h2ueRxOxgwPsULSB0J7RbiXmkT8+hRsymw
gOHK/UIZSIa2SOfAdI0prqh/iKF56JTrbfXENYCWcf9P6zyMybuRfN8FJq1Pj8Y3ZPsa2Kze2QN4
f32NlGOdTmw724DUUjv0j0gHqImQ+LRhR5sT0cXYyMBh08sKOkNb8OEEQjA3DIFGd/AOoV59cwFk
QUZeYOdHg0VOQ55KdaVebXLP0aMvzZqev5zpogCW99xYcPMZiEi4M1LLUbtcoAa1upRZyhJcANjs
HQkKSIiSUdZ6egjTZso3jEbURs2pP81KVKjofJhc03PchIQuGems5OLEnj4G0O1WaibaQ9ZiJe+Y
lLEG4+bYiRwn/6o6ziMuXXgDfiRHwZoODbHTp9uiRGycp9ah1pv2cCHX1T5mkRq8kKCucki4Zd9/
8bEhdDMvrhAr9yqBv0V1BJ0PsAqxzBC/scpG/rAyr/h/1PHVfCcJpTMNEuSktIa5q1oHKL7myA9E
0XlcaETjyl0I/r7+hham4hpg5FRfLYStEgSw/vM7FOYY9J7Ru1Z75QRR8YcuCclosMDgDHPVpYcv
lkOT+8M+7sBntgc6HxVEt1Rm5bv2Xn9cxwochKG7dp6zhoD0OEnn/fwYKMJNSzv3r2VtMNDrMBlE
093sHob4HMcIupIpUhLVfyGuL4so8nH5v9PN/mqyjouC79KdJ3OM8TaBCNwyco06zP1h3FEgPceU
HuO+o8RTanfoJNrbZfzqy19fVnZkQvy8Nbo6FK2pTNev++3FmicT9Sw4WHVCoBJr3WEqYSCryFCH
vcuha4J+XQZ+uYTj/VqY9cQ84NkjXi0ztiqDmdLjSIeswKWX2fjcYuYauEdMO21BD4hwHjk2vz3N
IxxsROEKFf6TBuu3xtZB+wXxhsUYkz8birJlYWZgbMUlu7b36ldbxHx9nczQm/ZByDDmoiIxIUA2
4H7IkjmNwYSfSisWodaW5D7v55cqLgWcr2/qM7Hsru5U+B432HnNsCykzFQ370z00J+74LeUoble
8DJcpGy3TSyxAT5bt+GZU3ChpiF+ojWx3XuujSAknCVlRjnCiR007DJKqKG1Xkt9s5ZMAZEaEGHK
hBM3fiWFpgq6es3dTGaFrJuGaCD7HPtplostIiJZdlQqFdNqMP/FZ3sJJI32a77z/+cRxvYTMttH
u0pGoZWSfZZNx5helWzQ1OfOSTYHZFgTW7jmMKIEhOkDuHYWD3/7AMHKB3vCDUEXg80D8ZX/JmW/
pZ7QDJCyvd5xps41B8RGKSsShZ3JIm12Nsdv3SJ6iQrALSFj1kd+fxpL2MRJgRkJqPaZ14d5wwPd
RB174CBX/U/jxFTR7m+eJgzS1JXCVHSTzHRsCwoujH3hROZOFwLuh+/wSKHD2W1azGHeHY9jBo0x
Mp25ikHRunHPchrGNkTulR5kAvoxyidfwjfsyhjp6XHg/ds3lGRkMxpVwoXmaOYQV+wgE9XhBARj
fm+8cr+IUgONVdS31p+Y/xwde5AblW1kNHCfltST67xY41Oi0kLGjpWc5w22fPF7jCmUJ5gBg7F9
FA93OJ4z/5C06AzkFs3BQ9t7L485vAwCAo5mtXULq3c3HOM6SzOgMInTTyRjJzhF/Q2YnmE1idGC
H3paAUPMJBtIfqUZVXIBZq6Jygu3J1Hgw/4jbvX9FGeCiVETDs+DSXOtCoDKeQqonBby34u5qUm7
lKGk8Ku96pA336uX3mwnZwdKzccmLMTpz2mNbCK5zUDhnbPbC6hHXQkw+1GahQif8HYRIGcXOXOR
4BnfRJVz6DPfc8YFEcLehEMxaLCLzGIMzDoZM5BpH6Tl3IOPlxYUzXAMy+h+GDEjw7kGxH9x/Cj/
TJAyI2gwPefWBJhhISJDF74UCSqpU89MFz+FDMJFN1DRkOe0ldHPsLQ2kIPieTW+syJEgkkjQ/HR
z7o58I33kc/TSUVssywppVYoElKZhhnHy8TTUOV5EVScjbcMMI3G0yOEGuvyTlpVdG6s9ScLh7f4
UicKbJnbGieFPK7FxcKABug6ddPYpAp12zPo4iAgwqT+3erlKDgYM2h1jtLNzJ/O4Ab9Zj4qIeUV
cDVQH9Y+EVcA1daTHsaRkzRT583jtUgGxFEZn4rd4MxgvfFy1tOEe8SuIvhXhPcubVLa9cZTpgFd
ZaXlKXhrIm/al0iYmWTydsB5ILZc8ODApfy2bFfiM1pu/n2MRn7wKqFEdJCf5krAuZ2oMvj4spV1
Y0F4ASc/V/xSnE+RRypkXBKriRKzB2aQC6wgPplJOg48bmVr6ovAraOcjoGyTQpKvB1ISHMv8RhW
XwKO9aUqg/IvoOwEwUMMrjqxgZV6s8ZV6srG86s6M8KEyCTXqUHkU6D2/FraF/FDb63CG2gwx6VU
hFKXVRaMtiFtXYGzsmFLDgSrhH4rDAXGccJcH6kC2Zv/Nn8bsyv8cSu7Lf0y2sBHLWUesOrn6SlN
mrGKN75fi2J3CPNQf/mJUyX9dBnbZCuReWFpRryEX90s+D77tLTVGncUOvjcthyp+2524a/FER/F
3Nu8Rp5KJx6Kpl15TbzEDe+OY32C8olgIYVP2AbNnwjcE4NKbvzuSS3dXQasadKLzwTF9rcMLq6F
vN2nZ38AreTrJHE98RCagZ4IgLmhpzKZwVC2otxw0fcBQ2DJeNXre2k7bJaIpbD+0qhuRhfPeeQC
hfe6wLgbhsoSVza3qFBljWt/JNxT2PiIoHnwCYs3YOIAzyzPWFtkSGccU6ZVtC30RS8JnZavyNHB
CAQGbqn2LXYSz/eKEQI2VFQ/YPPOIJAxHkbAH9G+BfJYF6BiuHO6NYx+tpC94MCjEfCgsEjY1CFs
zMwNaaLPesq/tlQdyaAIWFuXdui+4iKDQ4W7jqIRly7PfPkzA3GhKgXypiDmEyf+URgkemm1XqFA
KKNY2Drvjy5wCIwmApAGo/EtfYl9pYciqcnR2gpYJGp64XoOtsxeVMISWtcd4hzpceCKAWeND/CA
QHwrz4EDztWgT9MgmbNt91PPGI7jipQwrL+U6a33osAMxMzYuzIFrVKdHIDp8cpaslXkqBY0SiWK
USQLqnXQlltZ0aaLDSdgA6kv18hJWHjc9oQWr/UFtEmVtnGQ+AiYKUYSj8rR59ZjlCTsJes7AHiz
TxIqwBX1eRgDlNuwYmuz6MfziOA6nTgFsnw18xSdlGzQXh1iKQ4xuJ512ZZXkv9AJnNkTOI4G9vN
DIEIBGVQ5/oa8AQF689AJ9E5UshZBYpyv+8LzHysV0E/EgiELJMq0zO0tpojT39TtTnvjF+EIXkI
z7F7L74Ha4RCpQWZpHSV+mDINFaHlhR4c7d/DEEUL97yF1zXf5aRWfAssIL5Vdy+gBAS22fuV/xf
xaycLRg2dK53w8TtcGeOMfi7VOdsTIc/tTxNIck2DNz8x/YMnC2pnnigiCqbdvYXJUtixVm6a9sq
23EtFQ+hYA3QYMRbSk6GClWOcGtuslxqAiV9rAdN452r6T6YqN14Z6oojuj5gzaejatJw4IK8opG
QeLyJB4vGYH7FAhj2JMo7rpblrChGlZ6gAaQjIOrFO94rJibltrHSoBEVFmKjjki6XCypPtQbevn
YW2ofkMd6ORvdhIMHoJUNtADOpLEHahlYDRWQ1Lvau3iQW2Xsknkk2YcFaZ15mqEPTv+L6TneDJE
eJaanSRja+iXl3WV4mLN9KI4APlIcalOGU+/DKaqhaQTNUb3UpIorHk8hrhTQJUEfvpyIAf+4SYJ
SZaU61lh3hN1+dcz5wcj+9+xINyHM3ewwiaJBGPigViBBEE6V0rFjxU0YFIsYSIO3aRh+JZSgXm+
AQpauZTtRC6LVCajyrgyS8D4cKpFsDVG6MjLXtMo1qwKAVsNlFq4PCj8I+HReT35jLDp0zIYtQdm
vDrbMfvd8MnjUET6qFXJBEAJUYoxGkzqRRX93SNzZpnTcKPbY7UD4RjoodYnWynplN1GEYpSeZBd
Xyt3ToOSTUurKnKI8/3+ZK9qStE+Fpz5MfUNzf7/QNR/EYukgx35sCJ7u4qZKvuu92ekaOysnp5Y
jOdguQUh9BCjxOFw40Rd2y6vdInfIcGU4p7DpGKgvd+wjoMliyo9TaI9+5OLJJPwGFFhftq4XQYD
LvIbLyEKM7RmTsU7cMLuKoyUvePy2va/rjpRxGU8zGsAn5eNxOhv+80mpPSit07K6TU3VCA1puWK
+FXRxuNBWDu8jujDx8NBCqKWCec+U+3yuVFnXEDy1rDIOWmTJTGoVfWXOA24FCp5cxEAJkLR6Kyr
T/UB1C/CrrimrnrMmdCClBXNv+7SUSmPEhrZPGC8IHE6/nbpfyhvHfWksnry0DyzUk0IgU3ENAMM
CnimC8OVy7tvFNyCLoOccJPm87WY7rxkx1s26B8gos8mlDa7gCxkFI5dxOvWc/IW7cfXNnbQQLLy
/LQfxdnmvGZ4/XEa6WJLGFYKoPOO+Dlr1JIf6dNM1A5cEY06wCy2WiLrGK5MYfLv+go0mVfLI0Ik
3lbXfwItR2b2hcbupS6//JDfA+iFsGUrSFxIcKKCVWJY9OZCytWwQivh65+3OzmRsm6XvrWaXU2C
s1Bx9zr41BEYyukr6wER6Jm3oXDzmtMn+gdyBDm3K4n5YCoee5f7DCno5G8VHJkS6py4Q8BGB6ob
7CAkKGs6tlwxjqkTg07GKGL+Y0sGg1iccC83eB7b8tKMixNuQIwWkiNXAPdxKCGHGKbqOFto1hXz
6y9xlYMT9L3uu5Rr6hTFBwCVwqCCLqc7bzbrWaZwcrkZyrHThaTt9QmlpZuRMzUyUpR2hzqfLs1b
1k1LS/sU0cFylOs50BXMyS5rr9hbf3up4kKxgyGr9B4/u61AIjcgG8WKjZXm0cHvQvJwUAtF+olL
itsFAN6eD2PEvNS13dMr0W9S/+uk99becRMhaidaZP8cP4SgC65l/cNNTfSqPFRtnnCphqHvPWPK
Jts9xOWkmEcBtzCq4pFmhEaqcT/Y7FlZTj2jjaC8+cFWLz1hUUzdVFVZ2H8x5c1FOYiPVC/p2gnm
AhNRutN7iCWZODCjj0i1rlNx6DTL6Mp58gnIANzCqIz/clf4LbSSoXJ9E6Ibb1R8PXsFShZEhx0o
Skt3bwXyIMFstpXIPhlK1KKRk15hKOzjgT0bBgUFkTNKKOAsZyb+aSqZlJi9PJObqOd5cI9v3sgg
VPlOyMJ4eeb7Lalm75Zz85yP67PpmBww6nOPZ5ZfvP/QbtngjmVNHlc9k5gFTOd6lY1IJYlgc0GL
gQbEFPdEvWP5FpueQkF6GPj9Y/WfLAYxbfkWLr1NBRIWj+8Iyi6dliHrbyo/3XTXyiidcJOCkb1K
M50AXDfFUoffdEyj9LL1KOlEdWpuE657yj9DfpqVnTc9wPKCggKufuVDdXXKH3UaD0kJebIcCZ7c
am6EqklhF6MqmVHNYmV77D/u3NQd+OvNuBSo6gayQCYU50gS4Qqxe7YmOAfOgc2sJ25KhNlfaKLw
TgPF6TphDYJ6o2oCOZE8mS5UHM9DUPMFeDN4cefonkFrQ4LrSWbTiStac6nCc5jqU+AZi5IRUz4X
3O4qE7ZLaAzKAS9GX0NNaycun9slmXSRgP9WGiE7JONgLIVG8d0KKWKI/5weNEcF46fyxRy4/HQf
na9lBnPF5LN+YZNpSDOEzgXDC+R6pXc7FXhcf8iyRUYaYclbX78piN1mBDS75DhPb4gmeyLWxX+Y
25019r9PDadlspNboEOIM2OLyKJI1Y05WIOEq8pLIeSMSGi59p9ZcTMVMXhboW458YRMzlsVY1hS
R6Ut1AahaAZUZtmyysD5gMeeYu+HplP2LXmjRhSIGPV0PcoCiT0fY6AvpHwlbh131Cww5Ynkllpr
jDZB35Q17/FDprTKNy4m+DD06BfcJVgGqMdZauXelff730QTcxjevDEUQDVI0xLol8g/kNiHWU8H
CMYlPuGp1KMpRXTHsb0Mfeit7mC1f4/J6SpBrzy7CKWQ9/PhtD0cl1gTLaylw/t+3v3htIg+LFgV
2ogsYtzd8Sf4STyxcMIja5HE4+ncA6Q4qgwVCr/3pCWBJU6gFLFqbu/rbGCCY4AjG6Kc1d7hhggG
nyIeFufTDGdXAykZ4mRXNY0Lq/hTYmyhjf79pEmmP8rvfrLfyYQqefBhDHWtz+LAXshTonlGBnKZ
wN4sY229qjTPAC2iJOZfjNmIH0fGzyeN6IiX8sA49lqK6rOMH0LRlmR7pEk7059v2Qvc/MryKRFy
LUdFez5ntQ+X94X3qHe4WSbbvKRnAp/qhcId2TRny2lD3R6jHm2qqok3yruMYY1JD6DAv6/4DK/N
AFeYCeN7Qjp9/hhsaRrsgemo2vrpQ1ZBzZ2TwML3BUIHC4u80N8L3o4we7fAaeABinPoB4xNMxbN
05KuK4Q62qYPYA/sZeluc4TTaLxP8wJvCvZeDXp2TpvxsoASUrsLFIokzVIerrTaYrqBKJa6ewnL
35sR4TleRPPH7kNkOV9AWGg2wh0YohoxeGYrkFFmPM4mawdTm1YFl89NdSWCPDWQICXq4kK3Voi2
Vee/gPfdoL+mxWcfZMJ6ke8PEEvnvnkRb75oSoooNke52FqtLXTGS1L9ut0v5Rrq02nQ8wM8NdO/
RpSjQuL8l5ojn83fbGr6LhfLfVDEj1AKuD24fwXIxudW//Oc1m4mLybFSMYZ5ZE9V0pWO+Q65ka/
bbszTPR+8AyFsTgoQDDHuOai+yWxwBwQvPTQo+mabQaZ95GkgT08qeEntJvhQLcQ/6TZVX6YgjKA
tQAuSzQCRNx17L/PtTy8UOVfy/LY9YRHqPOJCIMtHEMbxnGLVk1nJCgJKh7/3Cfv1I9Opl9MPnwu
zM5JfW8kP4rhKOyNzeJ+MxdAbzBe0g4EyMrXYnY2tlH8kXsALQEi3ef7m6V/szoOagJemli+i7Cz
re6PmhnX8mQKEy0NUD/HLi9Dn1/eNKLGOJdXire5sbXzciujlkWKVxjNj178eGq63ILLdtLJ1nsi
KRQEu85XzIyMMYmK0eqpSfprTM1PgyRA87+z076s/7WBAF4qGGka6iezYoewdCDBnsTJhSP8tkpN
xdLl9YBCfhix3PY0cLOci2nE0DEbYUQkYseNn3sJjCSRJCXnlIRCcu8CccSAKTsI5a/xmbSw+vjm
VH026NqZYB4tnn66yNinMGbvNVF0gF+0AY2nfuPrhRWNio5zLAFSSoMQtv3wvuVo9OkkF9ZZjMs0
lz4VlkTeGUHSBvGxQJbkRT/U3ZXWfjMbfZzdQlJEpjwRO8N+6ML0rAVTHXLMW+7DdhlmgM3CXsI3
VcRpX+ryjgDzkmlMRBfmmpmbvAbpWIEWAuS50q8iG6hUXhNeEozZ0PGdy7ZPkME4c94BYjDUne65
WG+Pu+67c3CwIowzklbrQhqHQaiMXdqFg9ggRb3ItUgnj+t2K2/6f8Efd8+3DvTxJsSCFHp4WYT4
VRWmwaTj8jWwi3+E4IXQOpvDX3DdlrtrWE01FpRyhlt5pUshDiF9f+wcXpzbCnT1Vg9YNufPjXy4
z3Hp0SP03XflQnp7WV2nUxJPiJ98neyo/AG7pJkdxJxzx/8KaxynnzHbcw0+4amYQZ9Q/xZbbd2k
oTxUs9ZR3OJtjqcOwnDHHPMNTt2zog5wCVsQiJ6NVzPHEZo59PRjK9YVdAbSn8DU93D9GGYt/Tc6
QNHrAroHEXPlYcG7aiCC1G+Ystii5dxKBOrsmGvjNRX/e/cDvqJQ2l9D+z/k4lFP221Uq4saUybe
b5OHVsMTEkHTupo/9xA7dYmK3fFgO3Yf2DzfzQAEOXWsa5NihTpDiGs0qfpDPW1+oE5/nyB2IDRc
UcGV0BEipuVIvHYuf09dSmSyU8Cdv55b7YX6WmkAXh4EFwqQrm7rBBeLAlQAvwSUGjQWhU4FpbIO
h3Wb406prHzoJpeOG4fXQqQiRa1J3y9/aBTP6d0kx5WgYVoVDHS6xVD2WPSQYuvLgWKAcvPtAj9W
CLoNc88o4lrXMZO6zPQ8hhFLEiKE/+O45t21txhPfNnBLiV2LFx4oNu+jiCTaJkpszQnq6krQPeV
+6fqpXkFkRUkRlCVU0NrdtX7H8WUH4XD2HD1VCpkhSmoad9IQtH12PQlGiUKDFeq1aKhq/kY0+Zd
p6aoKr2OxHtPcyYAVVggNfWhdlEs/HAcuABhNlJLAdYJXSOG87MfqOGCjaNf5SkZi/ceBQ/royLH
DbKlO4dPr42qswE9YZxSz7XXJiY8v4oUFulK39EHG7tL+PrKNSbQGeUoSCYjCzTPheoW2vYQfd6X
MhFCx6tRHG9I8Ozz6pnl7Ds6Yslyp0TVh1KsLwDd9gQY5+moEYM4ErZ30AT+QkwAqyJm88fODbAg
QeKT/5SW9vSL8oz5k5LnjoXmAvRaJLqwutpmK5WkwzpoKaZvHm96y3Tm+Eeha9GCO+gGuQxIbPJj
k8Sqy6z5y/GvnkgzP/tjOntQzWsqTElHZ0uBM4iFylPc5ZclPF+F2IB8tYEGwBG5zmRTJQYTOJ2m
ivT6wD8qbBcvivSNymohOlM8UbgQCSw3hwOcVYjeT5oX/6IGqA28lZU0E+XvyeC5hk2W2RiC+O5S
gK/RGI97FlGJPFWLEuJp6Uan83cdlLArkynlul2PRyXFCoYtS8V3UAAqOk8GOoJRvIOls8TAlDHt
WNwtgyR6jVnGIuwdvX6yA1YiwRx31lxt7yoRoz6CjIQf7xTFoBULvbiet97yyCEjrUiQQra1BFRV
ifqKGUrSB5/dVqcy4Fst4KcU2QdJZk6b33Y/BgZ7+0Yt0eN9jwEAqUcDoBDoKhZwIXOlENfY//xK
n2YHVlRduId1P/ESi8WfgzyWenSwR+6eKE99me6MyyLoBAdCollbA4da85X/cS+AZfSg0HkkPXMp
6HCaBWhsESmAVL83AnvxesFvL7J6L+d4a1l6CmZKlOVB3Kt884/Ndpwyqla3JaSJsnO0K8pnGyKu
YOOrfB2d7Lej6RkkgxJVr2Yyr2kfngCBCWwAABgUg53CWx9XLpIisa0zMltPbaaveZi6tf/MDrWA
n7C1Gq8lQ9/lRA79g1q9sVLvzn3MS13d5+gKuurenvQJaF7t/m6wSIbcreqR8Fs2345BIshgrKYS
ZJEtyTNQjFeZbgaRD+X3LPo9/9E/Scg1hXeaajD3kasnkkFzIfphB1EqPLtA6OhIga9O2J335K+K
EiYZVdkkpjAaqLNXhU60/qU5qrPyhY6ite3EyYESV5RlpMJdBX4MAFuSLFVuy0ktqKrxHsLWmTLG
gi0j/ozCm/wx3+NO6+BFN7F5bHljjHWwkV/fA5r+FzitB12F82S5RgBjwChmwxT9T0WAUICxuTVL
mkqOEdd7l8t1Wt48X5USrY73KbBKWMB67rQcOmbNMw1zmPnCn+1458jxRs5Rgwj6G9MzizXcogG+
MViQipoH2P/KprlW6uxZNIR9UJ3wNfz4QREDfjReX9sCacTuCRd2LSzpJdNDlPki0MkzGeqnjbd4
wWjxvMZ0zGvgYyFqKIJnpbPhBmKY1TTxAygZSHmhubByKBXh/1u7ldpZbvHFXwxvbL915Ud+aFqQ
N4/FPdZLCHPH5n2I21zzrBwDtXK++tc1E6oEA8jJPpyrM/bOZcCmjBF2oMeiPCNEKyFR55bjBkoG
d1GPahY4pgDtCYo8mwKJrbzgRXnen3WaoFtGGhhkBLnsypsI9ly73tNGuozA4bSp62l/hApG2nDc
b+ebjiJWkXBneVT06OdyHyTUhjaSKQ3nay+E9Xu7IqN1OIlPidDdzS2wU+ni1kcd9/AMr7s4fKCP
WNuoFI8fJhEuTfSW/dGQ3rnc/qjt9sb1fpi7ZFmJ/hHdza5MqPVeYEQBhR1Ym3UeKFIpYVcwi33E
gNRNXpbPTRM7cTWXrV7eKnb3MBR2aiv17EMzCUuUh2nczYC6evLDzmUvVQvrX2HbTMu7llgZ9FDG
PIwXFruinpGS6CoBh1TMhXhars3/zEq9/4PQuVz6RavwJCyGATU0+QWv+99lHTSHgyrMGf6x/9Um
nVWug2kEQHprn8PJvJl5BzZT/Kz8COY/QWmhLzUS69n5hNaGPV0Dplb00ZOElQ/4J+t3V95PDaVI
1icMji5AGczDUKVlAmFsCoP/TXDm9UR9T14y10CWr0Cj0H154zw8rtjPc3FUqMK28LFQLxV3kgUr
o9Sk8gDNjNR5RcILvqXPQEg/htrw7ltZkP1f+IDQMxJTWBWPPFDwlERt3xGetPFzP1wv0LH9WWQd
17HLGSa/d1343i9VaminyUZaj+ILNAcYZPhhrEQLm6IpYMPSFmmeLFO7eR0QsyXR2zl8PhzxKhW0
trczptf9Rh6CRzSgRGO87ILknOm59S1TL0NDOTmYU1vG7LvR1H0IFiTwxRq2qHtDcpXWQ9MFQidm
Ie79NvfqsLcsBzu6AV8iZm7zj1e3DXX0WphxjQHwj+x37nSM5SJkLxc1o/yOmcXLpbqQ3VDQwqcP
1l+JOyU8822pBN+9LGGhf3mu3YTPSGMBw8P09FMv7jUWyLjIBQWXxu5NHuhWCnAOftVeOkdBLDRz
Gw0s+YtP45WQCiLfBxUo5ljrmG4KFxgUQg44b6hL/zqBJLkwkqXk8xn8kurMROvowlSpfeJ3/UA0
xhozkbfBgrEzng1yhCUtWKpDNLrd+AoXFO277lwT05uDm32stKfIWEx01MqYPPc0ffzAlO4T3OXX
mpIL6Dl4XfcEWcA4WdiK4AHdCAiZ9iAmSj61ZrbHVJdlAtHC70cG2hSvAtjSZyhF76q9Zmp7a1kP
31OLFdK9ziL5kpbPh73NsuBfEblJUpfVoUjo3GWLpow9uY6QjirgA2Bb9MbKszhi+Ne1FkRRFLac
UZf0Q7IDWwct++newx30uClIe+e2+Fwc3hp1Za39HTrL+XavER9GHAZdEIvY737eR2NHH8vmFYc0
NQV7fMHkw6T1pU856kD2O4LBJDGPy3C/0Pd04twCaV88QpZJUINNsWwLyPnmArJOBaUWqiGsEadW
4oLMReapPNpT4Tt9b6zYu2wRDNONFw5BbfDs/PoTwqkIDShupGOTWXWxllzFtADIQXimLoRsYM8Z
zPAUesWqXsoHKGFCpV23WeBZTsAK8WvThUAKARPL3Fl3n/IEJ+prSq7x4ZXr/3piKZnRxCMvZuXU
V6ufkI3XyDdTZwDzR/J5cXuPQcfwu8bePyv8IK56Ka1KZ6tjSHFPBHkU73pVWPGIHtk+fqWBKiLA
A7lrHaPJj+GWFGjUB51CnoGGlk+gb69NuVS2+jikXUwJXncmGJuWztytx3m3i++j2BVy7Vj1Q+UU
aiaIRyNrPjVAikNUJ8vlFFNdQ+sP5jbnP5rex5c54FeLYKAjx+eNlFn5LhJPrvre3ikVWardZnh4
M9kJymMMbNiXT6bWuv+c3z+64EEpahQVxsHHSc6peLUWoIrVr44WTz5uYYIx4aTy7lWaX4xYxMpi
EQ1MYbJnzXvykBHDPaVrqJ69UlRKvPuVswZWlnx1yFUX1TX0pQdWe0vQOc6FoZY6teFITqP6VpHr
semb5J3oo65ynu/NQSPkNkeikWz6DqchprdDBbpiK+D+Y1Ab88aLtMAkD4lacbnz+jzghY6hAsVd
lhKhDH3BlHS+3CChnbEf/MKJYvrnkVRsKPNctmRSYW2U7UChVRup4mN9hbZ4vm0HDxCnap91xm8p
KxG9aK1TkMWRqY62hKfOjoqokgApFxO3q6vbpSiaHVOV9tnNnXfoEErs6ZZy39NlFl0DXSFALAJA
VSQjFeRHzp3HbMIp+0eAMHwsjwD46oeEtq2Y3Siu4c8GG+I2HeOe9MpjktvkXya/FNMtHzNmoBra
sty9NeqPiASop6ytv5yePw4nUuH8hZw8DAsL79UWDe+yWoIRd/89O+uVig8WeB1BO8Zp3lx4J/KV
F6vcrSFkze0MqbsUPSIUFpPeoxiUK5CsH24jQrMnpUE9eq/Qr1rNISktfXqnSOYW8IXcE+NvvpBd
5m/vj7P017TmOiVHbyJlRBH+sjON5JWjfowqP1FsCjOqGcx6mRhnjTShngAExIzNh27kwU+JS3Z+
c9RV7M21fhAbkp2xz9nrSytyFaMvsDk/kThtl0wRytURwbmL8pbBCZNbmLxrpwb/WbX9SCBaYCWI
zpTN5IlUhLDfE40fO78gwqT/amXBhh9sWrzn0ITDIvwbmDRMnfZwfq57enuRNgoh18/WwdDeEyHN
YcJC1UbbAfWj/5YoIsmZAATp980GKg0QE3X2A377Yi7+B7Nnk0CIssXd2/zTFllpIa8RxwGRb7UN
PKzd+vN+sd+VFy4/ZweTIbQVIoDDN+65EPWLSuiyS783Sssz5B2vA5g8wHl99fSn8omIOjOyrKbV
TkVQzvYi07S55pfeZYgkKVJ5OaAikjWLXJXR6LVb1D/hPKOBSOsZqMmA2LEFMRirYx5NNAXCFI66
mY8T/LqhTHOxmqn2+yQAzZWPjf0zRBR/IsnVkCK9fqpp0UnBmWjWmca4p/spccphLRyW/m8T3I31
H5LpLtC1531nR88RkFgRjBY02sVqajYorPTRDDY2J8ohCt44yugl7LtjhoqIO/ioRYlzZZ/QVs/F
hF9p+j8wjSmnqznU2CBiwGepwJckYFsbOPQzASt4y79OLsSlTCmiJW8F90n8F8HICfoF7WYJZyDT
olBcwRpdFRjTTSQl3nvpX5XtTb2P4/HGIJ30hOTTn5PrN6sjAVFUMn9eilJM3D6cvIW5NkJrX0SW
/h+VIs7j0BfuS2KMZoz0D41FZonIWjKkqYSBuVyE09pf1jBpNuEivJt9z+7ypj0FYI/u5jOAReU6
VJT5UG90IxdkRK2VNFsyqGRkqHdmhcLJtG+XwqOhQ2OO3jcvKzzB3eJL/NIp8Ah63tQrug4/L9H6
B3y9qGOJkWsEoa1C3j3KJMNtov8Dugt65LXdKqIDRr9niDWiLL7Kzc6m8IFGppCxQJncOaPDTzHq
2HtdpPF0vBgqwzbtzZvu2aZPp6HozG89CnjjvQuPLcI2PqjsMtsl1a/0Onx+andnrTsyea8s6Ir+
jINDipsn9f0s9av1grvnFWquPb+u0jsX2hMgrE+21hIe4t+0xd/GzHAUzXHV6udYRfQcf6fFWaM4
Cu+EpKlXin1f5RguOEaklQ/8PIj13MhM4RVKXAUMWoNcAeiJVHUKp65xFtDXDznv2gUHN3GdecMw
+QnCMlAMnPjgmOF2x0Ep+rPvvg5OscZDsysUz1nOJ4Cz4DWH8kbJOQLUMT6EoJ9uRtej5GgjyR0u
X1G2cyU3rY5I8qFg2axUdK3KhrUcnL0vPLFrb9JOA1LhWm7a0pDRqyfFbqsi62doFLD2N/fIQ7fT
7hy2YZ+3tJmS+JjYoonL/oATMEGQ1wxVgLWY6cMbi4GSn34jUwrnNohrHA86Qc/mIl2dtmuwT/2O
tow2z4ICO0hUqg5mnW5j4vZTsYxIzlVxKli9NTVbkWRpEFcYjuxljr4f8iwLYUBZtrdetzWDi9Kj
uzZDSOVrmotQmH5iD2TWJKO9vXuzATCztKXYx+KGyNGszndT7kwCkFxBuYSPlJ9b6Lvx/6psUXLj
pnEu9+iLMa6nwHsonW0eYWMU6JHDK/ApF6PVfbkMWd34byTjCZHaNZbzhG7hQjcWJGyE4rDd1f3M
ZewtXfvzCaIR2fjxu042XCzoBYqbiE1iRtSZYwKXw2tpOuKtHHyY88HYDksluFfonKuiAxctrenR
iUSzXkKH2N8P8Lso1tyo4FFM4pQftSBXKpOFR22OP/WCYaQcusXvtHEn7OeUlSsfGUoAsXcg6ekY
bfXdvPlYkbgOSa3IkKxUx2mDMaWAggLEpwX2ZkcqrzYc1H5IzqSe+OETejmrqvAYQpoRoXRD+BCs
wTmFHpXzTnzskU3WezNy8fsHH7MYWp+Kb0Db2uKdh1710o7K1P/QiozEJU8ie677Wq55Az5Fi7cU
fTqsw1uYfA/xmRDi39JWDChUxJZndbsh1lDe2/PAFpSHz2FytUqRBzDFaTCMbWAQFGO+OPpsPAqr
tOTmD8SkyEmDn7PdGdhInG4v5CvGoApk9gVejex//7eMqF46CSd9lFGHcFydYThpAeTyZmJ1a17B
+5W543QPMmv41j3HjuiQ7tzjSdLvb/QqV43k/pN/QSudIxtTLr2ElBm80ghAR6JStJHFLM0NnmbN
k4ND6fuBV1rrzYtHuCo1QJib7uHhB06ld+FYK91rWyLuCS/A+8rWLsZgmgAqxgvOiRibqIadu0/w
pfCiPs+fyPfnWFvq3BYymnwmQajZLrYDvpMo7kxSqV3rqN8YDi788xVTR5xDUXW+BI4bgaDg+v3x
FyteyLpAOFY2kMNX6jwj4suQV9B4+/ZJFKAxzi7cK8IsAplH1uyOtLhrF2gAH36wK1v7VrQwBugJ
TIIgGBnCw9Q1NwrRu3dBEQLevQmQmor9udj/M0ToFK/NhXGJ7ibzr2MjSA666pOFG+rjHe1adiMS
70ZspaMmOC9BsvbdtNtCSxXGZYuP916TjITrVAr+U8EoH93xnExQ3R6+RAlF6BBErxoZxBOF+Lbi
ChJ+/+x/5Z581UmY+WRCtsyEK8IrHq3GNqbAPo6rP7oH3fQD/9zttk92jwmvyU224tLa7dv0kYhG
GAYybX+sjLfQL/fs73txe//HcgPP2D/cjyrZm/UQLZCQJu+Fnw8h1WceSU21LobKyJDtvFMEnJ4G
XJ+KVhIvDr9RG0U312Pe71U8gt9u+okZwIi2nn6OC6iqZj0JMcGvs9A+b7/ErZ3EJyq2zF0iUHrK
M5v6+4neF6CPycZcx5ERWt5zmJdXhgyykFtobcodvB1LNNVYyZT+WFSaBavk2LV9THswkOTifnMe
AuYhzozBj7DoPgIQOUBTUEEx8ckrXp3kjbzvLy1+FzJGUH+3wTGd738jRbbkd+VJNORZzeeKISlS
6cANJCIQk+uzsDljo34AFwyCzq+/y03YXXnORtdZZb48h23meH1pWsyrnKJcYD6ZiCFQLfzBUGX3
7QwJgSflxmmZRGIzYl4NTOKiZesd2ABnmd6EQ6xcsypdp2BRv6t6U98lUGjeEC4lV9s1kZBupb8Q
GuU+rasYhEkvP8TR92wcjCU5PGNaZQfEEhfzojuaELnlT+RZKJZdW0fU03yQ+R1eEokDqJaHKbHD
KhoiozDZKPj4INzDm97qucP9Zufwd449GP8IDWJdbtdpCStJS+MFik4DB1Rj+wUXTNx8lFbEOjxy
xCfyxluGNalxvKZQCUMQZLkv2EeAaebDPtFNahBuMOfljKLI/j53JMeqywcZw7LhOwCsmx56XIkt
LlRGUPh+KGeRHhWVb7+MUchBqr+halMa7GPiXyafKUbC62fgpriiAsy3pTXwXmseKSnw3mHeYkdS
V01fwvaBFoW2Tqy/1t39MPj9iEpplsTMIIj8Mlut4zSofg/iK+k6lnOWjkB3Y5EQz0Vg/9yrNJ5Z
tPvldzT0coMzJJjdsriFO4NA4AF1KlLFruEJXAnDvnMB9nSQDAvXG4tZs0rZjMcLJG8e/r5wSXC1
fI+u9Qx3rZmnJ9x5xWqM0jbPuNzA1dA5FEBzzI9GZ901EHhWApzSE9zRS8LPXtQilW/rdaWtQkgC
2JxZLOLWZKPr4xO8vWom8OYhDTXpCgLhK7s0Udc/xxtVwgo/S9Yzmi3BU4iG/QnIs3ETbQQkQQ+8
nYdl84EoL+E3uqukJ2yDIUDW1f4Tn+hsHkPh+DtWCJQrr6HUUgQZhKUaXqk6bXm1z16uXYexzJfa
f0e6qFkStUO/MsLJ6UBaXWKbH/PtF6qoRpMulBDAqPcigp48bI8YTZKewzL2KYk+EwHEBOKTRLMa
+Q7cDnKyqmcALAXnDDQsM/hkM1tNO/LWdvmh6q/ARYlCmgQMpU1lysClFmHtVqnbsscuGbX91QkQ
Jd15QblEoOW68/oYa2bB0DYAQIFEj67GaX4UV4QpBXbEhqSdMjH57Z3716Vi4GdlaKkBKFZwO7QY
KKupcSgqUCfOD/W9z1QV1b7zAOrpmmrXjYxn0rF5tu3Zl2ySW77e4Qrd8t8ts5aSD1eFKYGXafJC
lZ1VXRKCGqosWsejPf+Bi0wV2ajiXXqVB8KScblv0bVDGFtNuxKlLWYQwLEYdYe64daqFWMsJfAu
hBiHe0t/KjEZ+fvKgwZjSGRRY1R27nqocdMP+x/r3gzcoJjI4hcPgLVx6OvtlA2srCFzWh6vqorr
+YssL7FdpisEM5YqztZAxmvPg0pLeDgrI1UXPu7/qP1nJP3l5vpPh6SmfH2vIs+XHUGD+UuGRvMC
zBzItmotdzgUsMKNbJ3Jg6tG5aaLpHaoZOGUUPfzDzjPqL6IiA4ZFXpjs1j/hbT+nM+TdYTiyRuE
u+Cxnog987sh8UpLukzIky3IugvYt0QdOl04zwQ509gvAaGh8uSrajaSOXzhJ6hsenvPQcBqS7Qg
fCcq8KWqarXjndXY67Nvzq8W5/QGTNEL5AWN/0KsKA7hh7C2I0biNW6UYXA/DtJ61+Ex1aKNjB9K
NPIFQnzUH20lknx2dNxGFkxxUnkmkxQ4f6fsKDvKky9LVEJpfD2KkJkWIbhH/qM7B79qlrrmWR7X
PTZDac7OiKCB+DqLmNQnPGwdTFQeBsmv7J7uoSIcK7z0YnxHzMlsbDOeaGvmA5UgVdVwO1j3MOH/
ooASlWS7qBOrLgpl3MdfqbVj9wY7fH8bT3W0xS5RoZKFNzGq1Ktm3pCQ1THQ96bdWmQy9zFdxhLO
Qmmx9g5RtxxZL1vMaIPuRo28w97f8IMdXWvASliaUT18BLrWupsUiZbAe8Gw1nmD7C+HtX5m2D3/
P2kuS6CUCEn4FJ5KBYqVkoYYiy0NhebOueYdsgQste5ttF1QXJfyqrzj789BEukLmCYeeQx2WtkD
Ea0gMZBjXHEGchgfpYchM5IuHFBZR4BKPMag2gvITFDmJ70nZIn00vL19qMgmnbhyh0k58kfO14s
mb/swATQdOiBxE46l8TQz0Iyt+dybWJsM7sqD6TaVtjZ+CtGQaXngtI0tDyfWAnN7TYBGX1O56HM
6P4vnllSr1Xo5sTe0WtdKpRARiclGLHkydgDjBAYqcTeM/e7ezDHOz2x4dLq2/cvw0gWY6jiebfO
6TOxuuxHfyjWZV1aWa/Np32e8XcAlPLinmCWgb3ejM7wTDUGAuqOqdUtfy6UhJySUVqZXUxlC24v
YY/7DJfsKN/0UC72ER68DRScaStMUjgAdLGPHrW1D295UastvZXHN7vFSgaRrjYK98ujPb2C31PD
b9pTSmxKThYm2VMVMg05VWUTj+BHE9zP9dMyhznpd1LksI1/97+HLxH/U32s9fXakYv7IiGxjBm2
kCQXnKi6Fb0nauwQWNIo2Fy31rbUrs7jiJcr9KCBhbeT/6vn4e/LEBba0WKltVOo789MhAQe4i82
roikWHTxg1sn6yv2idcim2wsPXDas6xculdbMOcxFPka7vs1LaJgV+wnt5F3T0uqUmYOStdSmw/x
6C3lbNQNSAEAusWJAeO3v40BdicuS5VmyLRqsDITkyjS9ng/dNeE59HzEwcBXE2F9+wHXHZ4Ydmc
8wBWJxW0mJ691iPNoszj44qLg8h63wwMzcVlyjf0fBzlWRzuVNQO7PvFkV4xHgFJRs5qGePdtFrN
DGePav5I7l+PJO6mp3O8w6p9zWK//xm1XoG+wvM6TZuvLT/JSQkiYcuo4W3deJ/uNRkXKwvCxLkr
+lYZFmgXKvT50e9QkypBoXmkdwWXBg7ZYx2oy1/M37Yg4UhDS4mHgZVBj1ZbMoEh6fv+fXLTaNK2
Wxs5cnEueTfdpRGPF7eBDmwamOm/tZ3nsKfqnpICuco5poUX8djPkQFnzpyVINFax3P/tcMhj2OX
ZNe53eQH9Ar5UgUyFymrZ1ldaYwf9jB2YrbH4QxOWRCpOXDJNMxVDjNEY7ztsiE8gsXZMUPy27Bj
jD73KDrxBKa/vgCsd6rt9Snxy8otfPDFtIO+mjG5lEAfQVNkqI4QX0z3B79lgClxSaG6W46qiFKX
fBbfieReJOhxZW2DgMkOixAQqxZS92DITvbIUdMR9lGDlF/fhKV3V94Jyq8ugmVbslsaSE5kUgql
WZ8dd2/LkpvrxjP1LDyeJL9StLGCNHru+tyCQ6RxnPzDR8hdqP2v9IevGmcAigbmwKfPnZ3HdYq7
IzznX24jJ/uwyKc9KqdlvxMbTzhZZsba1NU/m3PeNYEOmcC6gddkGQTd3mRuX/ym86vrsA+bPi2G
wiKAHRWDfp5K8i56Y8xM7DhGTMbdsODP4/mzXL5DnWUMkRHI4fBzw6B5Vds9uKLlOqE1SnzTMdUR
7FOuqDfQvnauMnkPLs7vXyCV/t8c60j572YR1KhFJubTIUjOC5+ucs5HzaFYHwEGk/Elho1EScHJ
vjWA5MNlHnKIHXGXaVOCsdonYQBBdmhSJnSzPMpJO92Q+thsWsU2nLG/9EttdCitxIfUbv+Rdi83
Fg40PvDrvzUnDEJbL9tBG6QVdy2qNf9u3gqhTuhkgTPxa9+0lG1kI9vTSnkHyLpnFHMaSP0DOodq
3PIc9SosQkjW/xwy1TRI/BP1id5T3AAQhydw7cUUm6WgwCmF+Vi+giFDp5nF4pWT7FnaLAL4eDVd
HzNvFU/ntZfMjLTS/tNyVnfNHbsHMP8hwO1GhiJ41+R6TJwynHitU8sew4xrE3x5YvtadTZUd1nj
OH5YSuW4RmGzmMSEqgAs/xfiVFfWIdbR4vNsQR2DhWCckyolcM7IGGoIs7knnTLqn8iOAcjyeZsk
EGTwfd9rY5jMjI8A9P7PB3uEWPIy+dbWaFvvouKSTc2itVnXboF3RFTDOE9WnmC95gC7J7P2gQLv
E2VPdkVWCKa5jmNtri9xxgBMkpBKYA2USHWU4V+UPfF+KMUuu+X8YZB+uPFe95E8+ku0ny+7QNBq
pspOrUH3Ue0z6/9uJY7wNuaRBXNJgb/J43rvJGKj22J4iGxD1TgxiI/EzPVc/SOv8Xp3ASRypKRB
5tdnhT97nBGBU6tlABuxzTikEdpvdvcF1OOs+GHAQ4zTxAJhPvzD01hLPypcuaZHJyoQqzfpVaWz
0JTLfrWx5VSVuGt5hxL2Al1iqW/PZM0DZPeuI62LsNFg7FsrD3eu9/KacaYlB3wsPelV/iECklHM
D0PbOh39tVD6J8sD9gPFjScNPXOEFM8g2x8nUln5ux9/dhOM46yWlNEOmik8fFcoAZqFZBKnKtU6
rrpHwI+/2cqlxK1T/f0MGbPo+j+JXjNpARZHOD0YfSghcEMcepueNvnLVSno8XoQcA/309ojS/LL
V1hm7KBT8uF+8KfTGyqYbBW/Bv7luJN67iFWKhPR/EFIhY4EKJscR4/W26BucJyLO8bBouWqexBF
gQUdqBkjr+uxOfTDogXGI8lrDaCnAvkhvUW6UyaoR5R/3tdFLoo6iNln3IHovmhe/WHu7zhQDIhK
6qKvT0B8Nh/aOigjpPAMvDCoRbMVaRrkoZLwTdMyMyt4nHU6lzUYeJvk36ZYeJwXB+Pw5x+vEBI6
wVIo9N+9lE8MRuKTPAXmdGGgYVcN3IrrVg3dCXnl3Y8Y8M2Aleb4qgiNLnZDSVUZlUkMDsoV6KKw
IT/S0Xm+KhMG4KLJHgJl4yUD2qlWWl3VKoCLwKys/Hapg+k6EWWQwUyRziH1XT+gJ17EXsUyqAUc
A9FC0X7jtS7xMOeWqpCD3dIodLOxnSKloIL1wMP5qV2tcRRjniJG5yRbXfX253EC+ggZVBg3ONuT
CmsMy6iq96NWWgGquwUp8YkuBEMlY1tKE1LXMiunjUtIa2XLZrvJcQczVGKn+SuOro8YC2dJxTEE
BieJyLkKIcB9ZwGS6EfxGRL0o9EcLTSvSl09TT1m1DTtQjXznpPOpihdK6gjPfMbuWnM+dpxOam5
7YOqqges01v0kTdqHWX53EljJgRNLTSG7PupfOCA4jGOCF14ZqyPIIrlHOqhts+4WbA8jrjVNGaH
t03c5BfypScPWNamPucrUb8JeEx9noqLO7kX+dQRViEvXaduX3fCfj9dqsIyb9n+wKYPaZWKPznl
Q1BK0UBeaAVUWh3vBBWdVnDeyEe9yv9Zb6L5QLub0EEmEXXDkQLn0s7sl3m0Y2R8mbTopeXXYjaJ
V8ntIOoBSAbppFg3VGBikcoVPrDxOvEO+jO455iXCL24Z6ZtuiJ5Y4tAks/p2trxLSu/4cEyINI4
SjuXouy3u0YoDNUXUXnZdoZedV0fnMx0M0X/QpYoSSuT+E/nOhH5GqNw8yXJoONwRhtv/SGBPS82
VdGUqiaYdKmrL8/ni2vegi26yW2MJy5sxAR6mMGHtgnmc0pspkBK5fW0XEk+BvRo2VqLBcCGEa+C
FZfWBMWydtBBC5iIWgP0MmL2C2TQ2Mw4nmFCw+T9LawoIqpJY+MUriPOa2755e9XJX6t+JC1sWSJ
O2c4tV2ZbDf59vXOOoaRfiq0PEBf6qjeP6rGKPteYNjKP/w9c4nWMaB6SSmPReCzJLWr/QdIbeVX
innNHxdiQFow8Fdg38MRTwaU/lxT8NYZfJ7XCB+ctl5yo4muAkj2BKR9F2XYpCMT911uvpFe2GQw
ZirKXDilhBgZwmnSoV3O7MOrbmTk1I5mGc7R2O62kCYkbXHU8f2pJKxd6BaNi5okEnVFsmEamJGJ
wBkakKer3mkr0F+g91VY77Y4Vo9NLqGvidOXGt8aBBnOVeZoqUgqi4uXbIwoyRr3z1Z9EtowyRDD
uEZvc1gtOR8nBaIDfjd14qKkxOFeYkq68yMjchfrDZI7BRPmG2Dr85aYPPhP7JofmolSBPFQw1xd
Jkk/9Haa234KWeh/T8+z3XFSZawEvjAekt6BcW0O//q6nvsYHk8TUKq7rlOOth/WLFuNY1BAgV1s
fCDjbAS5TDRMCsYFbq42Uv9cSMvhOB0oLo2sMPRRz+UD+gm9bRGR2e+2BqBWlVlQ5q6K1D9piMJL
Gn4M+jlBclicmvxKax1Q/mmvF87IoSHBJDNhCtXEe7P/gw4Pth2DXItpwWbiI7WPp+lNvZGn1RyK
9W1JsEWH+3Mm59iXCM0LflkJhOBMiiPyD6TReMHmLVSbePWbM7dPxcW6qXomljVVl9JHxziqjMIj
3BlYkOqcsjkWwfF5StCoQcOtG103YsaOvmHOp0uNtFwVC/Et7UKPekn2qUIPAPwk7gA3S4uryRqM
KblERNydhPOb3qEmJodkn8TiQnNQo6Xy8OUMQDDJ4y8NZKKxIVDoC+YnILt1zWUOtkvEQMe/lOvv
wBqK4A9j5HywknoCGbkQlMP32JhUfMNC2ORDIRL+KMWVyyYAsN03nv4nwqIl5doecWZL8VjUfu7H
m8PGr97+Za3C+/VuObLAXmS/YcRqwXUPNsPMXxjYmDZ2tlsic/JOG5sOX+AKk9IBMhOLXq6Ryoj5
Xsu1FnFWoDj2jyxRNt8rfbslwG/G96dIy75g/69w+2hw3c0NHkPGHayJnR7/OlEEUeSghwgb5W/n
o+T7w0oqggJxdLnwSa8lQKZUYvJJ+TlMOOojI9vGze5jwT6olv/WDei6maivXvzycvl++uqs2vSo
mv+sHgVNPvUx/AApU8rBb2bFtCszLnNLc2qu9rvbFkovQb30LUwJhFGe6oGSckDGEamE3DST9WS0
SjaCvnXwXjyQGIISlAGTBzLo7mUqrfPK2l9mlva+TNcRGVHd6vnXkTlStdGz+CoBwkf2/Ly64zo8
CMIVDpP0HOgKmt3SIym5ZYS5dlMwYVpvlNShjL3eSqwB8cqkBMv1mxTeg1oJw41vl6f5Mu+3cQ3m
1J8PlZ32g5J5IdoCbOBm+44WNdjKuHws03QjojSP3PnOMuncwi2OcKywTrDHHzVoo8dhT8rjXMC3
h+4pLD9b+UQqaG2hkCAj8o4fi7Xml0aFdZvUGfEqPgz3eElvtnpVkwmMuW5dLtEDY/0pjn3flniu
P8ukjHNdzh01SgxCdog7CKaAiqXqygB0Z1A7aJv9OCg4TEeZF6BhoNAPhsYVNxHpgFl96vBemJZg
uJJdmMaDLARE8mxjNJ5Y9GE0hX5Lfamh1E4jfeg9ooeyRimyaW4nWQifKXJnuE+zZsM8viDdZ7MV
qa0TvMNoaLBAvFwQlq8HwtrUxdJf5ePkb1VGbJKjjOTNfYj1iI/tWHfjdCyg2nRg0BAPJMFBZ9EX
p7+mEdm11FCy5CF2vzfxqhg4pa9t+Y9Z6oYsG4UMRhzpHr2JAMxC6Q4yBCbdazIRrj6SRNTQtjKo
6dMiwyCYaKywjVX+niewu5nmD5OXXhtZRBzBMecM3nV41/cHj6EKLgHrv54w35xO9QrpR9DK8NhD
Jw4iF7YHtVnyfOcWhAWBcEaMyTLIj+gVAwrq/IqqhOJfDAQzwCicaEVJx2gIJumK+0+iboSoGM//
V/GsVAIP/LcearP2H/bGDlGEvNws2ZxakMCNY+4NmdmwIOj75iyD3lF0Jc1hfNvSaTcarU0G3Z+c
1o3YY9wBSekcY6TjjbpvanJJJgVI4xLAbnlajGfPTcNn4SV8FcFwyDG7Iw3kYYIcwK03OostXwpN
kD0PiPKH7Odaks4D6hpX15tWJW05awcn1tc+IcbiRR/Yy3jXR0zW2KUAZydGJL9MM7n5pvdKiSNb
B19pP38k8Yeph0oS3zkYlDUksRHmtC38+iEOLOxsVQ6I96WxO48AwyLbwziNxeNgEnNvnq+/rKKc
BOZAVGxIQzSfPMO9hVi1xt2rqtf+atkILHjARonz/W8fJyCqeCB4Ls8TwZ9WeOAxwgA3IIrvwjdl
4SGnI0jvmetWFHvMrslOeMLC/BZVIJDxaXoK22ObVJ31dov9G7ZWnQuOmzl0G97ZaqwyU/Eszq1y
Ck54GurKMN0RAMAzcmU/syJAisBzGR5xyfIuVcYgNDaZtxY8g+dnuvd2c/jKYERS2/l2cM26F724
uIAkQZXZ30TmNprWYPQCDOughAiW2BZbyS9ceOfyjAsNnKTlkzj6VSqvaorCh/QAyHkyIZywzzFG
g7Ez0j3BZY2UmmsygBn89XmaNqmaaSYK1uozPIZZM7D4O4snoCrmzn0E0IDPckz2VBJ8HIt8Zw+7
K+a3AVPHEnqmY4nskFdOF/uK1iZE1TXmB/rod6LDmIthH1QpXs3jd36zdm5bGNIW3g5oDRF/zzkr
oxDxKwSyebrWEolvM+um4RXcpt2Ps/BV2Nex1YYdr6Z9r+GvrZdily6oix95FOPR8QWGhYZ9OZnv
dNp7fLT6hRTO6F3kmz7pE1OxnSQEBZvBnfiWB1ubSQqtaK8mVtvqoJO44YW4W2ehvZl/jk7HSu2I
6D/EovyrSb6AdpALS+UW83EtBZ4/ppqzMdBS9Y1FddYAXfxTzMPIURC/pq2ToJO76B1lHtHPmcs6
H2jPNV/5x/UCVQPKCcJ3+bPMQzxNzuaI9Du0DzQSQRAVxj17Z95T+VAL3YnjI3TB2JNbH3BAed2U
Adk2k1X2KlXDGfYspwmWnS92ADMhsG8707+6GTXn3rpwLekthKMgRQkBOeUD3CzgrQvkb4C7HHgq
vEzM78vrzCJ3awJtMbTcvDv+mF/pKR/BAUHfOt24MPzjuijQU7BGoxZZLLla1ZjP7rBN7rPhvZwg
PmNuZKUxEAPT/p68oP7YdGNIMssA7H+YYdlbBdlAG/Q29gGsE7U5Pi4nSTHRC2vUXA2tPO9cLaAF
aZVa6gSxXwfntUyjB6l0iOv0FLUPXfUF2kNbiXBLr+QvTrY7VUQ88tBVIgd0IhGu/WiKyVU58EcC
qQSYCxRB7cjWiulaQebxd9bUj00yWf7iaoBk4E9w3Se++cp1gZ64D9Jm5WQyPHx4sxmVlX1Mn6RL
PT6+l7+bIkAtv5M26fWe3kJKF6ub80U4lfP2swZPEXHvDBjDpVIJNE3iT7p+k1Y375awK6pwWsRC
XA0xozLhQp0MZr+lXL1aTzQw2OB32efCY5eOxZf/qONWYkWXHI9Zik/zh5h28Fuoh78VnpZs55+i
lXEPAMB9sThzy//Ch4O33LqtvZhpxxR8fMeA00SjGz5KGQXsyBd6md9PMHVfAhR+hI80xNzaeAhR
dcb+v5lmARKYpBTucA7yQtLD9HS77ZfM8DWpgDsQtHoI402j5Bgt8NKb0JOU1nS2e+DAreGtsJbM
JNqfruCTJF0BKD3fGhFNPaZTMB5PHva0lfIi7n5VnYRGL0tVAiqA4K3SIq1Dl/RyG4OGJawdbr3O
Do9g2d9jeH63FT22ksqaXL/sg7DtEQ1e98gvq54dCGx/9kv6/POiKQkoosOqWxZd5Z9/fCxM9Y+e
odXgXnyGp0hjetdYY9KX1QxrDKQal3TfWeR33a8r3pDFrxyRYmtwWgaS3BNQQI44eRPzC8vY6uXV
IDLBJFMXgAV144qcvxYx2U06peUfolBlQ5193L02j6R34ufsNhyZFWtEjDWc4RH026PtB9oxRvEC
U6I8wAX9oSosy7GvCR7soTIi9U//xplxEHLvbkZiMIftwh9kmf2jhH7J2mh2HVu/NosAGRbsPmF6
o8x+Zo6y64+Tem569KjNu+Yo+nPxlcoOP9hk/eh+D+960mqGD7j6trktNcAFRuRuwOrRrAgyLNoD
Ifo46IglI1St6Bbd3l/9CNKfxL33+aS9jeb7q6bloG57H1+9Vg3WBVA0pVXDJ7kKg1276tPdF5vL
fJAr2jyhUTdij7oLV/qDookvUf5pRKVKZbWAX222+dbQvjeMKWJGSkYRkWIS5omsCvlN1LHnz7UY
SO1cgxQ8grA459mgig621i/olCOPNzV23Xly7wUWrUG8voCAHBwsErcuj2dQUTvXrhe5T+TGqQr/
1DKhiwtwu8gDmFXKHTl8RAesxBtuxYreIGgDsXkxABDRzBz6lIEniEq+OZzC9TJMHkKrRPVjB02W
Avorr8lEuRwpe3ozfflRkx8UXL5wcGaIaES+koovUA191KyWCMUvnWOkS0CKfICKHo7CQbo2NKk+
YgUe0K/O9jebBYcuPLTRaALFNG0/2Xseihq9feiaN0pqxuf47iiCVdO3+yIhnbJ7awaIoJLe0P3Q
1GT23cqzCvyacxy5qvJ1fuBsgkPMU3jO4QMWFpIhtnp6JgvSKWlAQAHfqcmYMo8ukZ4hOmhHWqeu
Ce7ZsH9DcDZ4m/WvMXavw4LNg1o37KC0lF3DDUvSsEhWiiE28SuSpmNySfzsSBCp5fmaT+Fwe5bN
gsHrBz/6f8Is+9AhfK6TBTE8uiZOXoKoqdYQa0hZk7lZRdYkvMSWgY59jNnCaxYSlSMI3nQiQze+
LZS5pOKSBh76jSheFaa4X1Av1DwsYXUaUW0yC79B61/HkUyQ4jF6D9pzWWO9u2Ya1WaKppzAIfNS
QXUl7OnUPZQdaQsi1qThUdo21iE4zYXhOVVme/GM/ru4ElsfJW7JYVGVGci7LjDWUHZWPan+uC3y
iu7jEm8jYRDOvL+fNsldZw12l9xSZ2l0Jx1eT73fQ+qRx3+62Mght0g1Ikc6SJ33BruO9sJ2DZIQ
kGVOEu0NB63/qHzuHekKf9CyX1q0bHqv5xiDact7lu2nFvP1v3ub70EWwPDEIUDUuetuGosKzRm/
ylhS41MAtxcSb/ORfmKsjg5gavzvKSifhi0QIZJ+PbGaw7p/3AvFkbBNA691WeFttK86AEamMufk
t8IhbGqrcI25SS/rr1Ba5jiyrdVaR7INIQijelvEGfiQ1RyJg4hvWpKxZqnd/g8y1ELcHXvYdo0r
i0kR87o+SEqj0MIK3huBLDiRXuskfWOV4IHskZ0ECcQnsjBQZFglt9ZP1sXtsjsYKyrzi8dDjTYh
CedMkOkUkiRnFvGo/eHcoH6XuJC5oKdkyR7JYaaONqObzYeOFUVTs58YbugfXp4RBE+gLdd5ftYa
pA9w7fDOPcxj/MEgxNBSenZhgtqrhV0l+lIM9HNOysrr7b1rM0riTuhBy4LtH+TjatBHzNiIhDJT
FvTHej4cV/XeSd+Is3rBI+wNMJ0d1FNJL29EsXjYJY61fEAhDKFvzsm18mOgvWHsUF7+RdHhV3xP
WwrNqdlWA971Gkub8yUwQN916lFcpwVeS0AcDxcibcVBrG7RTcjBBW1IsoUL+/6NjbLtTNaex7QF
qQvCAt93qiKt3e4kfst00/pt2MSOuhY/9Qr1yeA1MAiIQZDtaj/dB16dtvqeKvKu+EdLLAILsma8
aBpXpvrjspKAbfZYIMXwgHrV+pQz+R+sWPAxJdC/wkR4Ktk6QYFGVnKpJ/kHqij4b2Xo9qgr/Sps
41a8KUJie3t6Srbe9T+RJF2aGFkD1GwWyN6qHzL+16j089tZ9PQuyAOlHfMJY7fwAlqGl1GjGdy0
gidbNfd4NK69CNZv4bkYnVolncIccIg8Bo5B9/cS8zS14J2AQxWaRXaASdydLf3ug7HURh/6EpUP
W4SKWGfBqqEgJekxKXLa0IwtpWFf5IjHZfa2fuZP83NxRtnwTmqo+3MJd6fdYZPltDfRZs8aBhgJ
GD+iqKLYJLSdxdSOwz40cb44tlJ1SUKpO0NRj9ZM0VLegksgdPUmG5g/eDKOCOvH1tBCJECbiFa8
106xGZawLZhuDH8B+g6FRITeBvNZqUMLZPj1oRNaA3HwpeK6uOUPonW4gYofGz52HB2lhVAtTh0g
GqDn/B4Q3P7Ye0zPOXoFGZaJCDpeP6PYu1zBED3PFiO2qgMD2gIsT8YiWnhb694JC8O6zfSmjIn5
XCSFD8MwLcXYlKdmaA6pzqLngUgtVVF+5VKSI5PRNf9wnklAscUG8vstrPT1SDmJEfO3/DUB3MqY
38SDkc6k0b1CnvesDKAouGVjMmaW9VfdhY49kIoc1/gmMuW+qacJtc4qfzX6bx+7F//ca1zbIj7m
3r8PqRHc4QRn+HJSZcyWO+RenW/nn5OV79Cd8yLWMefPNBwbJ1nObkAyxezjJFOnfPHa83TJtxgF
zxagxdiBTlc05smFPfvjnlvuC1gyR0sGi+ULGF7s0EE3w4s1FsMoRNLt3y7D5PjKNS3JJ++l9f3q
Mn8Fof1D4CPjrIN9NwWZK+LPelCYfolMha8Dhf2EE9izBbO0Nl5jqIMorCwVWBPpIEj+tklxBv0N
SXQb6FoLhF1sFaXZz3v5nNM0H1LBQaUaOvazLAGR8sxfpGaXkaVJvSZt5UJhRe0OBB2+0kVWZi/J
lJDg0XNUvk7T7kQpYK0MgE+UNjQ31sjPUbj/CQ0bCwH1B2egYcX5+GBwFcIjjXScrWIKC8iAr+6C
VJsTw1nMPZfSkTfuQGAhbCex8oldSoKwvzNjee1kB9p1oigclueXT18ZCo1sHA/JVGI+Vu0npcPy
DXfVyAEA7dpP1wr22lCyXmC3KBJ/5w9kThowgaKddJiS7kS3mDvnLsXuS8xsF0CLdmtFQrrSH+61
cCwPJ9xHoXFm9lWxgEygJfW0j10IsEAQh5rmhO9QgaWE/9vUfkWwDaUzNbdWSIfUHVpnW4AjXbTK
zKbpf22BGTTKaL9EeNnq5d+qQ2/9fOjcoW1/pNtcpregAXoJ5ugc46rnsYL4g9OKh+y3KAkIwRpC
wCQL2j0OAfT6phjwiozZVYgS5lsckXivGgZiS3l/Ux8iBGxVqZ27PH89C0BNycpC3WZz0/ayXYKx
PmvRN0XU2p+2qRdjK77Xw1FTHNCBSdiLFZJwcR6EVmzmwZedGiRaviGCL0vC/Xjgo0sgoS1ufSX/
gxhd3Ztrqvg1DrysQlAb3kUY9Twt4Ds6juHcj8s1kL86y1Sle5FxwNH7dGS+a1Sas80HAv+FFKZe
/4q3JjccXD6f+uk1n07WwznkVEm+P59GMDSLCYPTzRgQ+OURH5Ke0jo1B01ymdUQbyWJPqljoToh
OjExn1yfTbfexFk4O0NvcJwhY/lO03golGEids3TgNSZ73Qi+r3m4z3wETpoH8zqj4jFmz1XUc/F
sv320iToLk33k1lU7cR2kaqaaakRpG+NhxJkpWWpBRCnYFnFk0ApJsSkZObSlGKFuwkeCFHuMRzl
jYv9vOsXWC8C68qVV1LT8+ahC4AZSEgRMWixDR9L2X4Kck1c76xqGjoc/F3j/rveK64HAsuF+YVw
/oGkGoJ0fYulL1dUnzBo2cyWGM0yMLxQvvyJjAs9UjvMQ0IQwicbk2RMrGbPl+a6/Ebp4FSy1C7N
s2GByJ6RNYpTtk52LYvlOLVa9YYRNWiEvyu1UfOeY9j25eWEidDMCaIzfnLT+ZJYdGDJqst54vmP
Fg8m4Le5vmYXJ03VOJLYVrjtV1N/Q+S+1EqWXFaYMj0kihchU6OPCljRyE3WuTmMlXNsqrkE5fNv
K/pyQ+wF0M2ldLFErlO4VxgemM6tE85+i9ktDCbGnFrrCszASjqAk1ULmXPnYMSkbuFOZQw3XJeQ
eU+wl23bnkTmrGF2NpDdZiiabIcWYX/cGvo3x4tHlByGrZCmTJxRFOLPyCrtGukJ9gDTRhgksock
i6jUzOgKuAHnjrQv3E/MlWJBaE1QhlEMYxSflAM20TCtvtfcmSw47hDf8DuC7Vl9YnfDSFhj+dml
A2BJGv0Aa5REOhS+X/AlDGJ9CegorVAO/U6tcdJFKNKuUVzbiR34NmBAz/Z0UBcpz4KiDt0kE/Su
U/3tA/LhbY4oMmCVlGscODog+kZozQnkgyDHOs26Xmm6tZU57emmUyWm010LOEYbuiu6qqvZZitv
ItYBNiPRKrYLHU9Jqh8meAIrSSbob+5/wQziyJxq1TeFHHhMxosmjVYmfOgKZb+7j6PyoX3qPkdo
oFwCa8jgSEWtIHya7Xsaf+zb6wGqpqSGOz3/Dp0L/ayZZZs3M9TDvh+/Ds5KBDWXBR8vDmRNMZmu
eKJqrUx5LmVNC3s60+hmUzD3P38dOJMjzsNyRvCsR5F8WVpq22qN0BueIj2OqAFZkcyh2lOznF6p
RIWs8vCf3U4BiAc134f7mOtKNTIkwIU9JCEx7qUi05TRrZYXEU3MYU8VwoXpZbnqCMJZbyhTJDTu
UMlqUcVWjgw2k7lhj66ezPX9gsGEvMt6u6Q+fuv54bT6B14umseahcILzqPk1cAaIbS/WXQJl8aA
CxfPt5ekbH/ZjPzoKFncbZnFnR2kkO1iXSZl5ivumEVVk7Xh3Vl58F84aAGm5mM0fCzPQ47B485c
PP/uUagyyTaisWCijO2W8bvz+PyrOVCpEdmn+U4roCriR3FjpPNgsCM8axTz9CknHHyQRVdaaw8Q
sYgPccaKDKEu95mpH/fVciuhzuAnN3VBN7XHSysyEqJzJ/aFFWpOhxUajiO/uhDstYAg/lIhOp3+
zryWPYZRd6gczVOqZvLVZMZFHjDV8tYTMBQD8nBmyY0CMygtkfsKaVNNcjtGgIHotSx1DYVfk3ba
Gao8z7o90I0WqqvGzVMUTMKeA75ZZ62rFkK2HYzzqIw4OihS1k+Cwmy7IL58Y+C3CqUjdUEuzBg1
FMNfSvy8kNqaCxoQrau7Z4W7LA0zHJIoQSSzWel+yOt1iqa2yadsut/1iYhVz0//hvm1SuO36Bmz
tiBNgXMCDFw4PdJ18UuPXYPdd9BBfuzKCSWNGBz6maYmYZYw7OtncufetILX294Uyj+FEHSXwQHq
/dO1N7clr96IS+A6HdEbdL24e3ut+juAF5JRv0eTgFFzVFZKuwsAJGgb+8ngh5yoq0Tx38/zj9Z3
Ve3Fhnvw8uUV3YWxI24Nkx0tym8yLdDsz8hdM/DWWMg91ycFzrXldXzorQQTVceQcNUnQVrNSrAb
L02rZ6yPPBuhlx4S8cOtHqF00yB+melaX5i1p6azHTGYd57lyxIgLGh52DJltsaYaRMUB/yewxjw
7cCjJiL+s/1DERukuBZ7ACFHA+VMjxYuoHkTdg8qdThl7VRYOIbbFYHIPKtZbHhBeSTLoslgoNTR
4eN87W8P2wuTioBHIig5zNyWwjmReW4hUEi3FbHlygt6EmB7qEwpYrrAe3MXaX8EXZSxwRi9vcw1
NmflB8yhOT2JuzDiIX25LeZFWHyqCbvB5Cu+nlGzDuNxYtJCUG9fDS7tIEqsgaQCIQ89Qq9s7Mvc
ooDwaJZN84kOP4aLyDrdPCn8LN5VclDnk68RYzXcdv4hM7DGzJg55eUlbd1aj5/nhW9T3s+RHVle
kBz3UFSg71dFiDXr/N5dpqGnehVZHyan/HHZFGYZ/q7CVkphvieycfgosRk0tOiCQmt3pl8yNx9a
nVAQM6OJrejIPu7dI12HeUJuUXeqzyIaex3gxDV18zIfR2qOLAHRvuDsEvYjgWv5FMnAGZZ07gi3
41tBGeFrr6aABsBcZVRkwzH/wBE1pBYELtqvLA4UThG4QS8W9WiCXmXicAMSGzAIaYEfghYcGKLv
dpGc7pMJUZxiErLPpmXC+nkte8QgLMk1+Cl/K5KyjQkiOLJP0z+xLIVbD1vvDjBlJ2vFQNJfb//s
8IBJ6Ypw3R+OxRbwz3Tor0BK7RgpayHAwMy6Nwns7KDgwB9G1oHfsgPn+zUmXVVpc397ZVoQv40A
g7um9g34VU0sUnkHgyZYE7Olms7xVkYG2Ka8iadFTv6u212QlqEQyD2uFI7Ot+R4wE8kxw4Mm9ig
3dT0maJgVu1ElKrj7GYjZm6Mxc/6gqGDZM3xDrnt8q2WHqWlu8DpjjLF/tnunu6kwxDPEFLoHHnh
GwnWyQW4KjHj3JpMre6Mx6TXX/f6SHQpObTVAht1spPj9ohRT5Ox7lS6jH62CCXwcOP1H6vyhW6z
OIctGLQmBO5f45C6YcCHahBlSHtKBCjbPlpAocKTwqB//ToQs6maUlARM4A6l8P3O1v2MAAow+7+
eD7G8wCsm+N7Ewb0yh9jfYoqXAGKdHfuiw/OzqwmzIwBXepRRYvzA4YsLmOF1sVcZlIWaAfdd924
cNPEuz4gQG11J4BCgZUM1NevgKD3QTJ3l3PVeGOOdu4nP0QrfWbqjB33EJV+xyCNg5zF9SwIyVlE
hihpl/rhhGSSe4zIKoE2wK0uC6O0194v127NhuBTYjkTZd/uMMvf9s1cE7gyaqotsKp9WiTi7buH
BhwSQA+CNRFsazgXttVFS8XqhvUVA0wQMnvRnSsMrMfqeBOl+XFHhi0IjTWRG7SDKlWJ0i46gYUg
nzIBXjstBgptUn5ynsnOK4DOZg7I9e02G7zSk46gpXQjQHhSSDAynwBFVCy1KcpgbKNF6WkxxMgk
CHVXMGLhnlv/v3NGSxLrKItnftRDbn9527IXM6aL7AeRFXJFEVfzlKiq79LhoOcgTQQUQ823OxhJ
QUIJmGqU7/04/+LVRAkd9cu7NXhyUxA1Km1BAZp9yzzu9gYfgFngQWzHP0Yr/UpwzA3AA0fqQQcq
WgQ8MmEsj4w5hBIFof7HjAoe5MKuL/pYTz/8J5sMTvHnZDFclDrAXEC6fWUtzguz3NHefjm0+5t5
YD5cTFKJl09+k+ClfQPiwPDT7FxwwiZISx6uIt9HIhury+AmQ95uiWgzsCR7E6KyYetA0/NxHkfA
wOWWYA+++yqp1flAtbtSg6IYxCkz7gqgIP6E/BPtk8cVnh5B2gteWVd4lGUcSL7RS+swqtD5GqD7
hJ7S+Lsi8uolQ1V3qO3SqOOwYX2pm7+z3iXwEkKbp/+039KOyD0ZQTtoz4hFTwgvDGBS2unW+uuf
DrtUmgGe5cIXL5h/A7swlbXKjKyAlQaNoXllt+kFDuZMr4VsEzMBzGYjw0W2EzM03li0ZSRJ6pfI
NsAtpLHTAsK469+qKw6lUI+Cxr6Me3ot2TKTCxkfh7ybPQPu5MWs5B1fS2RmB+kNWHIpSQSHU/02
qUpaNfSZANWv8lQcOykeYoy6ZxKTMUsyeSbkdZi4NEhS3DnH6AWVa2aPk0uHh7Lm/wmp5b4BB1xZ
6tT3+Ms6oiatrUF3Dck1AzusLRojapYzqfQCr59VRIdwwvK2j4emBMH04st9yWtrq89tqfFS2P2k
L/f+JDhRo0Db7ErRWGPJEe7y/J0eMoxT7s+SH4/Wj6Eo+6H1nSucQ7502JY1ZKcys6PMFaVwTBeV
z7+ZRMR608j2kdA+KP+V3Exbvfbc3CfIYVsNQ44gcMNa2l3A8pw4RuHKw3PJROqMMgiKX7+EcAnK
pm1k3U8LnzZVAvN6B0MfF3s13RrWMtkWUwGGUbteaeZc7shKMcByeEYlJF7+vtBC5cf7rZ6XI3+f
Zz7qzKNumjtF5zNfm00mPiiE7dTVsmTg4/ss1ffEMyBVWTdV1NI8d/TleHEWU7Mwd1IqRHM4Q/V1
hjRs1q6bD4xmVn5ub3hAjuEQc+H32O1GUCRUpzQtQoEHH5k04Etz/RSYx6OLIJ3ArYGFa7Dl52nw
NxjzSpLDySBMKJuoPvXCKctMRLG9MgqzBQ8Fdu7dWstTDSEpMv0TAtMgpN3dN65wiQOnLt45a6sZ
AWDIjHSBdMcN+6iXO1w/7maIB01KupmvV3gdYjhSMg5+wrAODzzeaRVEIjyerRkcnCUxJ+LGXuDt
ioQt3/JQeg4OfpnJwAHAjWCNz/3l96wAzryPHai12Lg1w0eGjp9eK/gJyc1dufOrdymv551ShzYi
iW5IYWk66MYFMKlsBdEqL8PSNdZ+a7NSqvF+ehfwN8olPbE5yRjXhA5qZ2Ws75Lwwl0kHdt+jsJS
misylUllHAPVt3XiCXMeydQqwZS47+FfTkmpr9ruDvInEaG8rra6F6qOhO3UrZzdJqyEyPA4aP+B
v95GYWPrI5xcCTXTQ3YHexY7EKpmDSLbzz8V23Z2yw3Wd89xN8+R9LWVPAzNsALiIDrDCJ8rMyYD
KMk2i6ihhb4vQ0bIgJ3IPcCFlhNfICeEiYKG0mnt5J4dFT2ZXgBcG4KbC9A3NgFWMb6dJKaZtiwF
p2tJGEW6YG9jcVXVrT2XNEd0gwsD50Yd5mKvEyQTw+P9gr8L1RD6EYF2KwNelQX/YnnsafSYOvJe
0VuRT4lLv+oqE7jX3TtCee4keKeokPq2P/C3Td0ABEN7Cq2fALANu3W7ImTYd9g7GoaU9HzqMv2i
5LNuQZStVurqyhnAQ8TwttqviGvWoGmomxHyu9uWzGBShJUo2dr5JAqYa+TwveuoLUae7wswDEcz
/ncNmVfitI12mkoBVF44lIGzH1F5J8ML+RI5e2QU3dOh4zEvUt99r5Ah7UrCIOJ4dZyvJQKMtXmi
67IeW9pkxpFWA/QyhRE6c3zDiywjdz2dp/H30G44gFErSHZXcMKBlQGKrAeUXKdQqlTlaQYXy9m4
Qyw4bWrywaDfHLOVjX74Nmi9qR+3Rew4E/KpnvV7lWegkjtmIVx6gHr/cAYxhTmUzPWvD5028YRu
wGg7vc5FioMtjbaMCKRQZyqIDPalos9zNKPY0dTiKptwo99g83BHToNY8T4EjydilpyR4hFP3mQU
wy2/+tl5OhQubw4LcKrQoiesM0Z45XuQwlTjzL5tXANos5G/biFcz0/u1ZL4FYR1JxPA+YPO+iXI
RPXTkku4CxcRwiqLsuz3L7jr6PRp+C1eFTRKA0E2w7YQqiCZ4xFcFH/ExH7mesWrbt+2k76J9Tqm
NdExMa+Mubp5170p4hbXd/uHpuXDFBTiqd8pj5hygAxEPtVRbBgNMFGy08kBWeocbuBelJAt9YOx
FIuqyyJ4rOZYSdL6nCdD5gVF7f9LHF25kCImrJO0Sy0JpBGlxxsU8v6YrB5tLSmEKkZURGoSoxlg
pGly8KaqaB79jI5fmoAfOyTZSPwxH5AhwokaBmO0CM5Iueae0C9zZHQ3b4HaAvZ5AVXjE+H2W72X
KqNL/ZYDK+WyEGIB5/moxZaHunL3tEsnSWr654xnzXVTjoHr1jKB76M7JOR6k+mNzwzUTeyWP0r9
hrKqEApGbLlhSxXMJ8ESIB3VFktXvX+NWNZH3h3ZgsSdGNmQUG+wNUymoL9mIzyuVm00eAv4akY8
n2OoHnolUhulWGaraEATZG9ICNSv0cWSLIPlRxef6Sc9UcavZio0nvcO7Q6Ry/fb/fiX80Ag2M/2
28K75ZLHKZjSJwlEG2jDFqVj6NefiJGph/7Zxa/lf/fnXFsoDf6/Y9EHgCbzMZePVguTSQEiWpWx
PNqa+I9EObDPXtZJfgDGqoy7mn0pH+rrscuwUQMRdUKu4cga/n+VE4shP3ES4AMyc+2ietOHzpR9
nQCHeJfj6C2c7IXIJ96ngcpaXhlVUqZWOX0Q20K9VealoJLO5Ov4iE2dX1HFhFjuE7KxBvHYcJpK
lvhxZy877mZ/9OrMvDb8wmCpymNhAYtsfp+ob3SiUC+csR9kwc80fiIW9kXAUI42KcsOx7rXb2KS
Svf314ps+0C/qtse06k7uoEkVBKOp3hQTqFMb0zauAkt3Tz2e6T5lEdVVUmIwgz3BVKjDIE+5dEi
YjeES5i24hMMEVaLkhD1WzY8w+STweTJnJXcwxTcwd1RkTn5/5geymYOr7uM5PTitF0jkZ+3uZtP
g4ZFYdceyABppIchba7mvchMkwWmoOlcA2/ufOB6a9K9iCeG+HuQ5upJF25PfDlIhSt9Z1/DSU31
OjuL6HYJKNJ6Oaa6dyC2Fv69CKXIxhZ40XX/iVTa8dB93IcP9IQOMIGX0p/C1L49Ejc22X53izXk
I+69vTmhZ7wuJ0rvA5XPIhiwHuPuC8B9aSiJCt8Ch8VPUA19fzB3jS9Lh2AeBDUo7SNprxrDh8vu
cV1+XEYvxrMTmIXRWL9BwvU+kEM8AhSsYLUMqOPN2xMIRQXrtqeug5wYm4TA+OzMUiGX8kGGw9DK
zsrbult5Ed/YOIzjnOIjU8Lw7AzEGK48QsZcprt8cb4Ib1lmJSOC3n35AvT5tOBnJyVwdu6QWHhK
ZJmzEvROCNuesWZTQuxxtA3yloDvOvTYwDJBpFFzOhsxvPGBRA1afeYs8xlzdSjTRZMdqLmYJ9We
3KoZQ58Xe7fyfsHUj3q2vosSb8JCTop2wrc4cJukNCphU6co+USooEHZ4/+5adxJ7I+1Xngdo0og
pMQumIsANdMKwbSomkXATfpGpnJvqI/1d2xeN0JcyQBYpyuq3R80uT56gWfpjrJnkhrZUthNBwKp
jyYKt+p6TQnAhF2DrcxPk7Bu8rDdEQjcp71GPtHXF0swBEkR+TFJ2Cs2aNgf+2t8MtD2ycJFllBu
NXUjqYg84y+4q7u41gE1U8Hn4sPQunun36eUfuweOKFKlztFR9vPtVFqLsEbrCEZGGhxSTBRVBG5
v/m7yj4E9J8k0Qhij/GGbzZHcHxcrfUq46kh41OneDF7/al/tS/fFD+/iA7vRbv/J3cOv3pjU4ey
duKDab71uGMWFi9N2UEtiVjFfZLh5UVOAnnF96PR8RX+QhA9p+0rn2eZ2hWBDkWmuChYy4zQPIUe
j4G5EPdcjr/0yR909PnFB16BBA+uDhkrkVldRTAAVtUkj3+EF7MdMx5bNN9cH+0etSIAo9UsMzsB
clDvgsWyf4JoEdSbN9ptXQ9yUupm3MzQyvszfVWiW4vsV7BjZanobe56NPJamDL/3OMBSq/ZaW0T
s6sxCXn+h2Pb9CwkKd47sPIG14FXWmF+2z8tvgisnBg0PisIlaqbmFjnXquJvrkweqH/uWZ48gwj
o2cd0rGZyrn3fV2qabYO0RDVjrjpkBimzPs1DOn36tpgTRkDGrAF8CEJW1BiIG/0VZpr63Sl59or
CnW/dzWiorxa0ZdtH8N1gnZUsUbg1lzT3y9wN8BBjv2HLukW1EPhujS4RlnhnbcD6dk6x27LZYCp
1GvAEXOfqw7X2w2ik4ObQ0f7di6b42gm4ZnmkzwmwyJ4HEstlNzzXxPwZ3tj2DrP50e5u6KDUOTm
4HUj276bWVpfrPBbCfCond/CUuvRPx0Zagd1h7QsaICFkj/5YvVA3cLTpktPYRHFDi/CPYTVFuxX
rVFxVdiZOacy6vEYk0CUX7wMd2l9BeeTtdlwRBgRmzhOC05wY/M//ecUq9hd6JWDK9N3m3yEhD4e
KFLwtJiAOSbc+pETpTzHD9ESo/cPJejGzwaC0+vIbNhkbq+Ktp2YQvBEESzbPiAxvXvmlBzrBU5B
ddZypBclYFUIStdqMGF7+bvbBlZ5QNhT4jhn+RiU+LOBeGT0GxcKO5ESVKy6njWTly3DIYM1VVVi
lFtapc3Gt0hcyV2pcC+zRPLQKqjCrldrJNAXYNva5p7xuuxnr/Rk30MJ8UBQ4qvz0OLZHiQGSeEE
fgB7UAWDZW6VLp+0n0hY7OrAhPlfRiarj+zx8hSdPCgs4Gw9JHvRmoO8c52xtygfLNVtPGZ943FN
jzNvqEy/O4Y15uBhct53Ccr+d3sM+FFO+rYLBYaSISwu2E8LknQT1H8TPVCh0PjaxPxy541PAeTu
THXWWnRrojs8ll6C6eUDvb8WsoekDet5YiMxHpAH3rtmITJpTNk1RNDPWkpPBX3hQ8wBvCmcF/g4
gRZpBnEI1lzA+bLxY1HqAMRKsBGzUllT8BOUJMa87GpQNUj+Jakwfbp5+5PHpz1gNHFCIrElIPe/
oh6cis/eCBmINryubXXJGb0gdvOHyMufbtVeTMuj5v9gDyN/FpCi5rI6WnXNGDlO2nXJpCKXzXOI
RDIXdBt1dDH3t7HBAt/VxaroxRfc/cHPv035jfmvYwP9Bs0GA3DShdyju4zoqLjtwblT4hq59pSH
xzAtSAIIvcO91oclnJ95tLY5m7Iijci8hpejK/sccp3v6vaFvXCQeAT2MuPXdMYAptHQEMSyygXc
9jUilmoRf//3ZA+6W+SMPsxbpzeGVZoKoONuYmaYgxmww780DL2PY/DJFi99pcRbbGPmB55jq2hT
KFgKjh9DFZTyzEHD0t1vjv5aYElm1T6tC6r88v9QyjWGk/6Qn5L9bHNfMfzBQguIvhMS2XmPXTFk
5iPyIjJ8v4ut9BA0ifTdj3JjNMJsfyW2dI0qwV22SGlTk/dUKxPJmAvz/9XvAD4F3njOS4shyMsO
KunWFU2yFeUhAct1XvfoeNYKXMsbVeYvBBfaIsedTPs1ylaZJ/AWVUe9tWwT/ApTw4rJWstHhim+
KBwnbAWgIxx4nBo3E3EGAttR/7nkEwbIt1zjuX+86VWIPYLKExh69q9A0kCIe4sfz+lJnkR0lN0D
wbdXO+KhIVRpinJbYRga0Yo14Cse39EnATrnDsdhFycH26SMa1k0H+wmtaWOl022sixFiUFkSwmO
ffiue6jCYFf/oTipXmqHbeSpDrlfDCAxQ3aoLJ4U9vJNd1IWpAxjOx9RVZcqx3bWUo4AGxrknM8t
+72nfX/BAsPEeANRO5xohDMDUcxTKn8vRq7Nwm8S0chXvuyJnhQJjng+52IbEJzB7L+AIgQG8+dz
vxV/dsGZoIMv4kYA/AK4P05Zqytqa2QP0D3x5fzYxbXA0L780A2QHSiyVQQpzkF1Kf78kTXVgfXL
ELQEgiUM2piWkelsRsXJWXp4k9y5vwMb0/sSD1cIq799Su1Qta+s9yDrmc3JyP0SF1cWb2+YE4sA
6Sj4X9aR8kUktwlHJpNGJi7aG5pMJWwtCfbNDsOx3KuRJRjmNtzHDrRn4k4OTbVrV/Qx4jTJk2OI
6NzUPLrBpbU0W4WGDm9Wydxr3EiFYbE+DOS+i0VYiOa3fNhqHcFq+8WkPoplfndqUjNVy5Rja+1d
pF9rKSCCa1swg2oj6IHoucg2tF7iDMbCJokd21szKckFcfyg9tU59auxkHIZn0XL23/V/nnOwfUy
dh8fd0kFDnXfFq2N99CLhpZ/jBZMHNkjt9XbAr5Ls+K+ROFDl3bM1H/hsJQqwLzuWTsr9ZhbkGDl
y+8le1f/sVlS3nDDC927UKyYsD9lPD3aPVlHtUVTW/Pfw9ZBYHGntyx8pOtqHYHlv0+YnekgpGii
cvKSuo32uk2P4mH4JJdGw7q01anIuKQTD0trgmW1Pp5k6hQ7z72ghxvX3e2nUtBvV1CuCvFI1QtF
YaOQ4OCMfo8/Fygk0pwfxflhE3uRSMRF6XGPK7HmjQ/K+3YS1sOIC8DqBElMVGVy1iN7O1Z0yZzq
edLbdINc0VXAD/MxaVsNLTGwsPu1kyh3yHSzSROIRTugP1F5TUTcxRv//og9AwDqKbNB1OtGZv/D
iLIUaYQMBpcxnBOkGBHrK5Dunjowye8exdfKV2nwNtU2jyqJGvtv2Oycplzc5ac12Vrtr4Xc5pYG
8m7CTW0RI1ZoCxSoessefDlxldkeNXZzBZlGKsAnSBcUBwMryGf9O9qM8Ov+A9eKNZsAELhl2usN
yNJZe5+xWz8eGMxN0VNe5sllm2tpDGqaERnTIOwSajIoV+wrpu2IF5Jzq7GnjpT72qX4qUTKXxeR
GJsnZm705e/Fm7d6Uzsgz4AjNsaw+M8JLqrGuxIFuzoTBTF08uTZ6F3PQKjfkS5v56QSvX7z8WdW
kcyC/GYwR7j3qUsPlCUmO/p7vO3k3rGWT+RezYqxd0tEBIqAfKr+Wm5ehDbOaJbrDZEQ/SFwDL+Z
bfBpVw1iWDvCMqCd8zEsitc9XDT558xbElwvbdFjbzVLiRokF6/koo/yx0Q32qPWEXzaYZgYHP0Z
+K+c7zs+T9piQw+HKgxD19YtX7UVGwNHh9ddsmFs4uuMIX9oWCb55yWe6yfy1u8Agrhqc6TB2XHW
Ua1EfmznRbW2sB6QMvPg4RWtGPPmizvjuOEanBY8D7QF0ID/WEgdISW8o6x27nh7lNZUlmJSN8jo
SRGWPRCNPQXPLS9KWFDdHJaCTz54ZDVoSEt5qUeXp608oUQenot+V109hzD+DZ3sqKokS/hqAOHa
C/oPuR33mlwJ/EIEHoABRk9rXyIqBmxD155NWagdcv3leOpwlJRipwGVBvZ9lv69ZurDvuxIlX/a
Vy4ukCFhReDuyyhWt5cE0Ajdijl+0Nb+OmECulQTUkHOYV9rWslrALoLQ5qSlztpA1YhM7bvWjn2
Nnq3Lo5nfrpzbDFOJ4wvvSHeK3PNK0VjupeQb60YNZ+bzzkyxsJuajgAXAoplCGA3DKkA8Ff8goR
QjLNKDJOEKqWadPHwuiT15QDO/FJfW3rmfjkMthAJPBXuJKPmX4dmmR4M1WI68aTcutGbSLVvxM8
DqEzQgj9ej6Z2S5DQSlo1N/uYUL16qGAPxs5hUslE7t5U+3QMYH8LGskQL863JRXhVqlVZBgzDxw
M3PrHrVa4rncu488wMEATxp6X39EuaBQpX8NsWWIfKuMdWKxItGdsNn0Q7lM7L4Zy4/P8o/JM352
2RVik0t2Sp0CV0NWZtgbWrCvjCouGqYItOXBah2sJ4+XrQxzfnjkc/Ir1oLQiPFNUiaq0MXweZo8
7ePawQHl/LHT0TetqtC05vrEVEzVoFsxhOQ2MXdmijrLDQWPVdVcVZLuREfuiDqlUCPwq0IN+h6f
VC3Qge4OQ8UOq6ql81a4kagE4HVQmAscQYtHV/B0zvxcp+c86RptJKc8D5dKCW7enodUqdzh9ut5
zMkMgu/vOPx/nuFoe7cPIMmAoffwCf2Vl8QqokAyXS/28ApkvpMot+2w28bu8TUrJI5zAj2+/xo7
k+ZTfZEHU2vjTgB7CPzYVa0G1IyCwqovoq/AW/aYBxVbQ5CGVvx6g9lVlOstQLsgB0NK1cwkRKY7
tXLHUxHl5HFazgDhARoaaTAbnvOhle/CtgL7oSHAKbbcaGFWF9wEpeEYBlraAbh/nlzoDHWyFkqw
hJRr3/YBH0w3k5m5A4NctXOuntz9GxOIFM8BX78rb9dwKmUcLkNQMJKccfU/nOQn/L6EMvDTPdmT
ow+i8PwoEgX28LNWS3qpWXPeJjEnm83L7xcDzm+TbYMlMUDVxbsN8f7c4mp4DjsvJzCJMjNh4PrU
ws0B3LmyEZ92XcmjEhFnGBPSrLTI/cCGUH8rM1bjZapD1pzVEeiDADpto+jhExK4UyE5grFGHDtU
OgohKAMhuDRW/0AC8JeCrOnJcnayrRdCz+fT5n1SuQVaDXMpBGmbpCPvdBf9Q1WBL5Pwl78cNBKc
RQF1551e4gxJ1/m0KkUszipiH/V4BT9vvaHyP4rZc2nbwNzFtGaPtK+OxqN8iYxU3EQykeOTZTG6
byjggEjthMv6++rAC1DndDKs9uQhaesQ//3HCdC8gZw+8muboQrT9nRRkpbQdgyRRZ0w828G45ke
Zxe7QU0oyp0mLHDwS36EJ+2n/rboMuNn7uCHMMvg5pbxyxkLVkGiRoFT4Y6plyr18VDiVvyjo1MR
X+HKI0hBED7rmw1vSc+YVdsCa6YUZLkyiRg5lM/Ve0BRXDuhBjcsDc+eCI+LBFsGEsMBHwfdPMAo
R3nMjQAgNr+cavDAb3t5xHmywlJfa/zj3WEJCPYA6EprV5ST9LO1sMo5hKr/xYlFDFnIOOShvgfZ
N/8QfkuBrKnFWGfVl9cY84VUJLDjr+LbaDUuCdNcw7T/KHfoff6GwRzK4xhoIGt2zVZcNelExqmE
zb9jZgH6J3qxFmjJuov6fN6mQy/Pa3iH++Xu8wr7/3QNrj+be1KLt/XoY/TukTMpoe6SVi57WKeq
6su7Pz7VcDGX7C6ViIsmM8g94gMSbMDiqEMV8siJTOtdhHgsI2sGgg4d0XNkoYLLbNky4rqSshVh
6AqHb/+D0JbcRyO2CAD0YU+lMD6345N7GtNeUPTl+40FoLTgSAhW5jRecz7TVWAQrdrmABF5e3X9
9a9R3jiH8WOTM6VV9et6qEdhdWd6/j8d/L4s7vPTau2Af3wFSsBASOTZNyNDLsZ9jWixcL47N4J8
vqSMkNQtp75cGk1jWwYdBmenTWbmZr/sL9L2GlSjjF6NUjNJLYkl4Ww6oDG3FA0QzAbOd3wmtAMm
1Pf1cvjrOBkrmEW/yIQe1BeE4TNyOVMalxx25WGcksW+1oe3ZRYbhlxnSQFTH1ZC3hrnPKMhhPq3
815Wmo3MX6Bjf98QNsqSZBJdBGgBbeBGTNa10sfG1cfD/5AOEuxCOfXmRv2NdKinBxrji5ZxP/yl
rObyLqYtf/tclrgfY2t2UqNdYehM9+bd1SPaL+zaND0D6bo4MA5YDTcGDqqB0l14moyff0URQMCa
iIFxVa/cgTYKs3K65PJS3WWtMhv8lWsXuqS5Y8w4Zp94pZZIWPay2NT1tQe+dDFqvTz3eqU38lb7
NWNDipgNyOY7irJkxMztEjxDcdhOHhgczak0xFioqJ4lB5VkXZWkdZQ7YUTfJ63kHfy2ii0VqQ0H
53tsSR/t07cZxbEKd5+36A+1J7Kp1Gi7lIS5ge62ZPggTukP8HF9KD2LajUDZH2NbLs6MMmTel4T
N05IfP5U4gg/5F0kC3xp+wiQXUWw56BDcWsi4o0zKda+qqy3a9fdz5hTnblUTClq2SbK2MGaP7du
rUSc/D3Wc6upFMhITKWFhr8jIDBXkh/O1uF0ZE3hLhfQMiyNRtyn4faMOzZ972/BfPkj5JptHcvd
Ch8Tf1rQdtce/K6pMO6pFKbIzxBmPAuaeRjpuXTZpu6f9oHyGIDYgUjrEimokTj0onQvoIeNPsCN
e6GdToWqx89VMInbNCnYZTWN3Wm8UsgCBIM4Xj+7Gvaetm8gWO8WUOZ+bC8PVyHPNHa7GarxcjHa
Sjlx1sSIj9eeS41sbUqF7bADo522UEXAxWczm2iV3ijD24kwIsb+9EBktTz460afUGbGTf1HzLVw
CJgHIo0Hlcx5Veda8jUnCUHtMKmc0en5N9JI45O3+HT84qpPZHMRx5IAc94Byci8CJuaeKzThCHV
pKBsbziyyr/htPfXXYGgLdqcsRzhinn9MvsdUleF/3ZmxLcc9KC1DlzlpHOr5JHCkK1xHGjukRj1
vSX65h9/cb41xO5Ke/j4OK7ECAaPq0qp6Jr73jLQ9kttq8ovbcN1mvnDp7vkeTgYyDiUn+UrSw47
154zCnCHl+T+ktU2bUNF7RyLNp+mCetD3d+i4L7/Lxg95DS9EtbreTevKM1Pz/qnNbr0NSubcjPj
m4Q2GiAyfke2weHf+V0qJKIaDFwJLnjxthto+hYY9vDQKhsqI31KyCdDsiR8fzPvEqYsWy9STZIT
H+RBNsM0hGuxaJGisiK8muz8SEbRs2ZDGNA2wPlclR1G1xFXODY8ilPuUPetm9goKnPyRu2mfnHw
iPA4iVTgmPAzkR8xWLWZW/4COKZeCY+PNNSpRpWNYL01KxQr17pSd6Gi0SPiopXszPegnRjZHLR3
Hro0Syw2P6zzUHckQZ0ZtJbb3c+VpIH8Bxsds6HWoeBTMNlOz1h25GJyiQbGX9pXCPjLRsTv06rL
zaTVaiWkLRWachRnVhSuCMIrbwVIDwZjQf1pGgyQekZKKkrLhfjNvjowVuxX6XM+cbMFfw53/uqN
yROc44JrWPfhwYq705LyNS0gNzqNCb1EoxXijUtmA0FdMrcUUwdRI74Vq/wT/PguxEdCdriSnt9X
1XeCCT67+/xcvRbAZuJFv5ntBRDWmk8eZ1Oba70PEk8cE3yyJ0u44ZZJDti50ETe3JJ/+yH6LNwK
7aIsS2IassHlaMihzl1jPeeyJWOrXS2ArBzW0K8ZyhkZk32p/M/MlcldS0yfKDfqPixhYwL0oADf
VqyvjZD/L+PoQ8Awc5t3v6RX5O3EQTa4dmR2/r/kcuDmt/1LfwsY37tK3QXisA6Sqg/y/QmmHOWk
Q8NtDzhNdfE3bQplG7H2mGjzm6e1KzXLtOGj1Lv2SuCb13jDGdgL3Ni2RffoaKagNhM81+dadvPD
t9XQtubJh9Y5tlb4rm5AyOEPM2V/Lf907ctSd2lbhV2RnOM5jjJTPD4j4OvQIX6qYRVDQTPkQxai
WLPshEcng1Lpq2Xy2BZrfE4wikCnyeRU+5llDZz5ZVFUu59kQrJPi1Cl7k90tfQ2UMethMAkqtuq
R15BWPm5vpmcV4z3/LssMABuK21mYmxyegXJMgo1zzPCFowk/tj046H51DdTTSZYhjtaD57teXXg
xgKEGP3n93LqzhtbgK1lbtudoZlFLa1olA+M/QUTAQ+L3uzSqgwsdwAtv1DpauWSSix32gbJAEK/
6esOp4S3s71Vkhf8PtJSo0fEYdU2y0cCOA7AU7DSdeSy463j1Z9FvkMR89wUrJsmryB/h0ipH23h
B8IQ4EuvHiV9hLH90sGGolIrnPmh7yfmIriE/XXsjBCG6RnALWJsFjt10cTJyuRR4pCEFd2+At1o
KXmmcinIx9X0pY21k/mjQoGj/2U7IHqdaoR0fsuASCDNMREtsBy0VYZniX70lqdd7ufoK8242ECI
piaz8x7fAYHL7aIOfxob0hYwnjrfVdUEMVbqCyNMB2VJb1E5xvRcV6GlMWqBZdgoc2gpD0k7wkYx
AASDZgJq6ghe8Q8nHQhUtI5RUpC2QpAHyTpwtpEbeuLCDN6gCr+1me2ayHqcYK5fpEeZ5LHGVHgb
ko1229AkAkvryL7iT/t36kYlkgiWkx8kmbzSuEmbu08fvwI7pjgoWBFvLTIYjBubVn9nS0pUq7qT
mqIMD7khUr+djzsPRULpD9TBIcuugG3IsjjI2e+tE3pGxxsvmXPGmLjIS5iUmXJLrY36HRwGWEtM
Wga1c73BnIoUJnGX9ZzFt0GLRzt43mkHfX3h7naarel6KtqdBo3GdYGKyqQrF/w8u5wSvfSQh1er
QgFsEjV8w0Uy/zx2WtnFwVkARHXSJDWOyRyytgG7onlLKTUjyTrfp+3Jit9QwDLXEln1NiTxcXTM
voTUQ2X3Blk8om7TJezgXpVs2HaIUN9gzqCX0lKn5hWHwctX53ah+tCsu+hzwvLEVEYSqWH6jyOf
0tsVMImNpmkLoSOHKnBTChQpPJlOr8/tE4OjWL2v9qeAkrxKPIlKJlmsKMfulAr5ZbhGSLXOkhge
ZeMbGhCkNAJBxPsMH9WH4gpkOg83r7TW54qOPyI3FFtCOHAb9hdSUd6DeHrZhI7nQYHAY4eoLFrT
oX7bDZrG+WU/VjMBIXXkpMJOCG/F32bg9uGM31eTffa5+fVIZBvoBYR6OggQspry49vEnAotQ0TR
tGqD6JXtZ9tMWHreSPT8GXTOvlZtvk7YCi5lgCHWGlRBFQUi05MUJ+khDHtXjjElw3LHQRope8ip
dx9vfJeGUvjrOjEGk93GqzI6mAm8hg0cMlGCv7Z/qkBf78wLoPcpaeQPzdXgtNs54WyQBD2jQfK+
A9f2vFAuHgDwP5AgUwPl6M8kYNH+XnG6ZxwOccGg8MjYst7VpryrEvasp1/oMXXzY68MyvSSz5nN
6CoQ8pyjiwmZ1NOwjRy3P0cRytVY5tkqsZkh6uo1SjJOjDRx8imYRPwK2z6luQKOfBiUno4c7crK
kNqw/cwFWFpoIIsPLgj5tWj4eRJGqx7kXADhqRegxzjiv+Q89GyhgrO2vBRoj8H/hLegaTomIc8D
uMGxSLZvkUZKdG+t3QG83erh901RjqO/bl5iUV78UADLRws4ttJHp8sLCnmcXhaOhWSrTqoA3J7w
P9kxZ6f9njc/iGtclmvOufM6oXGhJ8pSdpMMAknFIDs3eSEaZi8NZkkgwQwOZ6cySFTBNShQwm9O
C3YH00xgtuPzkzkefRgwiQRPQ5MZE58tF3AeDtVqn+jzBIK0Bi6bdf3Kw5qWdtAC8QOZTTMCNhk9
+Mc5wCO5/TzQ3BxRrBrst4RiWXmpDsOlfPYluxp8MQ6msg62E6/09kMypjk/I1SWFHUmKy/IrTma
4Sg/PVpVUFy+pyMh6h1YgywxeWiq8/0blRcn+VuOnmA8YmXtPEOXUrAFZ1xH1ER/Hfs1ixgTKAyY
JCYeGZBjJV5rydZ0EGjHqPzfKUPljBPckC6l56KRm4HuC3PqEhrYCxhwns5p6VatSwrLW1zUIvob
XRvYnFF5EmnKNEDfpdAR7Arx+fUMR1ZbtAu3fnapBIdz2leB2tA05hTf8dNev0VQu5JCgXl+Lr8G
hZDv1h9UkkNQS27pDipbqB92hkIip0vMLpAI29fSe9FFb4/K6I1g5p0PEDy/nLLVifPTbdoEImhF
1tmb7c+lHD/P61IG4Re8BMkaeXhwm1EoAsHGZyTvkCyuaLaen3VmZ0aw5RbNa4j4g591obHUuFmJ
iNoVvjaN9iYY5RMpRF4ymN8JLAxdII+IQU9w9WoqlG921BDPdGQ+4ZvHqWdBjVNzq+vQMqT+J9J4
0/9pyMdp009w5JvuwqeZDo7dU9Pek7Oea1/rzKf3ahLxU2IY2ndxbzFvkeXQvgWgzheja1whZxxK
VWqX/AXwFx8s9TEoUC3mzCtC2Lv+tUfdWfCUT1OmxvaNhmeAu2q3rcU8sb+bxlQBvPxuKpR1umNW
U/fBIBp7MBWj4hDFiZWM5omBlBte/WwjCjz+zq2m7j8WX0uVY5c/rsY0PPFiyV7b6Ijlrim7xUaK
3JIaFdrJmUtHutAZtL+Os8zOV5E0/bM3i1kAB3D6ZNbjklzLFNNz3oVWK7zz3C0eNlV8sYJaCln7
BCP9bKrchkknnvLHuE0jh4z0Bl4X4VEJQcKwe4X4lsKFU5X2MEG/Jw13WMhyAfZufQzKHwdHKCQ5
zNJmuJ/YRKUFDFBlrEQnUdV2xQBqCtpNTw2M56yRxtuZup12l/SVAw6wg/5sIRz0r8J/J5LbIfIZ
V3nKZcyrZ2H41Enzva+/Izgs/d1PBTz1zUzC1/DRma6f2IZ8ZHylWPq+Zj3BpIca+OC9KtAwxFBY
I37Tl2fn5sMWuxmSAisYAORlgpPlaufc+HK0aSXVEVcdDjnnBTwTJuNvSj8F/0LggmhAdkgivBYp
h0oMGR8WHfBzhOWA5VUNRHJRZBRPWC50z0NyDoguh4+Mwge1uDVIIH/2jupH9Hs2xeGg22z/XiuV
vpGXyNsZlJ0YHGLxGSttwa35TDPQaMe9AbBa/rg+SEVK1RMDb0hqv6GEWYeTFclyMPoJZl9vHcEb
ZT6fqjGX9epCeZSSqME/+HiRhvCZomZjLboVejY/lqXuJHUO4uUUfMpoaMpn4jue4HoiUA8+804i
S+B0AzaOOrDXIJvfpnBs46l9ydyFGjLSlyK6DCEV+4ZKRUeaLO5tyAkJ4blxsCncvSsazaOs/bD3
19HJerrTAKu0N6a3tjlzwXcH5w1nhLuCWfUT+ocOpFDfVmtf6AXCbESjoPblD5wqWUiHmNH4c845
EJP8XgEDhvRRFDgZXe0SSMZx8EB41Y71SdiyM5bzVZwDQ8LOn2w56WPSpC+fidrJ1vWvYZok9I2O
WKcdRUIvK0cDj0UBd8DLono8n05fjKps4Oz5vzc2OgyJRpAye7EkXv3kcYEqjWa9laPG1SXHu/lJ
jq9/FtHXQ89vzgjv+IQn50AM/G3u2ncUPmaU6jXibzmJoQOmWo5No4Z2BUqiaJAx0IrvOFyg1/+y
MrFWebfQaDf1UKdad6do/m9VHrT+evha4SsB0bOdj7rt1oqzlgQx8KEC3uwJc+rB1GJmfbyVVkoP
P2SxPXcsGA/F1tHir/P0vRjwjMhRWD87uLRsMb0Ul50t4fMx2TYKFCqzC1xvX4cBX/McfkNasUA5
z6r3fj+0rGaWZp1MSiyguo+7lWuzL0QMRBSGHT3vdAM8I5A+3ki0tr6n8mx+vKP4BvqL9VsWmA9n
yQN+oFCODdMx3yFYORuZX4mJ7UDh07LP7YRmNmkbqFNdtW/rIGbUBDeZn6FedGTkmr9B0katW5FU
vtJNUqEf5grJ5OmQaaRtYPf4byY1oCseS+ILDnZg/jQrAinDYtKJIq77I5JuWbVUmrvUDJzaT7Hr
ugRw62Bu+8ipTF7zRShPHPxtoUPAl3XbBmhrWUI6fn8jh8I4oj8aphDNHXseUrUfLO3kRSHlkVlQ
WIVP79WCthUndvB1xP12QL9WQzP+rubhhpoLa5Us22YiT1ohRTjvO/jMryv8ez1TtgeBMnR9Qzmh
vRsqDCAjFumWWXrXOAEsA2nCxS0fbE3ok3+1vzQCfvEIGXBbXIu9OxcuGxMij+MJ26CrXWWTpysi
NUS1NWyz+TTP+eWa9motxd9gQF910x2AzFnRHN8v0xTYJ2Yyaz8pgaV0KiYcDPhWboILjnYsI8FZ
WDfnq9moxGF0VCShubn1D+yNu2YOdT+JNa+a1+MP3dtqOnadA/B9I/sIAo65ln1OvnVWAEm9Z+H7
CQuRm/YT33iUMraLBYOpMXxz0HSaJwIkg1Q6vi2Xcsio5hPH8S4L7yE6MGKmuZjnt0cqCkQwZZoO
Rv4vP96jIL8KGZO2rX+mvlQ2XgrxdAgCgvBqy5wGq9t9RKqHzvUzkaTJRKLgRatu+WsOLrd/JCNW
9xeF52jM+QiMZCuWABs6BoepqNk3enz/chTG395L9rlPGpZY8ix9eUsmT1hVBABCPzV5tIJMZCFH
K+93CI05xYhwh4GlrSz+GYmFEGzmuSpUtHMojfyw2DQLBHWylRMuVnJQcFNq4WvZyLrJQqzbya+u
pECmCJwrS4C7jMz/I/sLVn00pnsYY4RZRKpPVJhK2hsHyZdGwR7HhCJ6VP0yrwZONh92ssr/6crl
fyi+TTfLG+WNNBIwepuk5lk+vCxKbLxpLpU797pgZzy6V4A5koY85H149gXLeevxy9ANPj02ZoSl
SKScUGsXiM0IYm33nUVcGdl4M/nluGWP95s3xuHULEA9TRNksdURQ01xS3ZHG/tLFl7lUecrDKIe
arlbl9Cv8HDehyP9MXERltX/7x/jsqWHWvOfZNc7ugU8q11eEtAVyAZMUjYM5bROgDxxPxO6PnIj
FOV9+vepZRUEhsTugporRm3KxwmvAMZh6VBMRJ9AQMK+RNOUh6qitjj42V3s05TN1+NZX0cDIjYD
ymYVLmFQ2ZnZptI8gV32Gv76vRbRhiedkGfw7c/I13zPyHekVBHgO0QDpJIcA1mDnTCIjdI6zOAZ
BdfRfPyCyChkTEHA3xDTzUcezMTIIOmn6pVAhHk4WZaWmk5Ef+LNNebciH+GlY72bcz54NElXWT5
4DaZraPV1ymNuKhPRBc9O4bc+nGfzMpDVUwa1Buhsj9K//6gOvPrEb96FWvFyYCvshA7C/9WAwwu
rETpcg6fDVlAZmMl+02RX5LTgzZtf1V+6Bk7aCSh6Xovh1df1RjCS7dIWFB5+BxUZUcMWQqJgjyk
QxhtDMmiI3h2u59bvfL7WQ2dQEohvOEfm2DAcP1Pw27HyFaSNaouQ/8nkWZ5/+rcPxFUpnm6ZmNS
4kR11cZzxaV2O+dmNQjPqD0TR9dgX9sBOVcSqbriiCrjLImUMz8MgI+G8/mHhPA0dvQUTmhlCHkr
G6Xa5+DV9fOQuF3Ge+omA8eBl+eaBAAfU2yDLAajaJnXB+B1P8QCvpXStHX0KzYoPFUxi9ScANqE
BZ8KwKjL358PRg4+MiK4Z0c9WSDvBGIOV1c9ZT/3J+fjW7Qqvlji9Vj5CvreRRLWazF0OejpiXZ2
FuKJzxWibKR1s8VF+FrhiR4R8ureRLmPK0lnCzued+rGmXO+z7o9Qvor5WIxTMhMaoysvbjGP3+Z
g52IaABMMh6pRlLqWLsS0uM2CzSWF303ZiMls+Omg+UgUkartH1SykmGBg7v5E+C4kIrT3j09gdd
mLAry6LN9/LgB9Z3GoQJFmRxdeL+SSXbyUtEhXlXp6k+BRTfYvoS1wmBgMtfK5WIQBFbrCT89JQ6
D7S3Jz+1Jw4xJXfo4ZOiJj4hCiuQ2+hZAcdYn5FLsiCVNe+bH7mMQ6qjfT6Pgx01Eh7IKqYT5/WC
uOguCw1T4pKC45M5WrOj+z0I0TPRjOLHRAAqUkNlpiilkmltRPZP4OUOcdXeHePYMXMHkcKJ9ZMA
R1mYw4nFC02qDvXHuFOjevATrRY8l+vbBVtGIiQxeu3czZLOkUGOy+a39CWnb01+jeZPmshGJvDP
TMpOTgpETC00ER9wgjPY1ISnvXy0hIIxnGltNWTcT+a79+BBDysaP5WGkMc1zhPT1JwQWWyyBSS1
b5nN5Wc3HiQ5riKEX4jv2BDZnX34K5j7D0X1zJ8+tFVnbKGMaYBRrFKvMCKKvd7kW4zTU399K+5O
PYu9FjfXbYnOVe2vIta8geIHo6vCnnR65QC7jbKmravGaUxC/oCP9duPw1Ir5Ham1vTAHpSEPAA/
cd6O6SevimD4V4XSYlJ4fxYebX2V7CKM1LWiye8ZVPcfxwwTDhgD0QnPcUVtZ27OSjmAdDfwoSIu
Bw4FqUr2DsgsStYS4T4qEMQHuolMIruPW5OnuYHXZ8/3S4WjMm4Xl49IW6pyu10Y6cKVXsr7wjk/
c01nU8psMQlrawe13Ts5f5T0w2Idcb0K3iSQwBO/YxJz3462pWhO6OpERXsdWlHwKshrMrDDrG78
Q+jXL+3TwvGb8MJS2qR1YFjDxqFkjqwj/qU+U1u9ZK17svv+TMqVeyUOd01wvW8KtyNc0RnM1sCg
YvQjUuGH+joEYVgrt4KZPftmN3LNsmKOju+0y9jsiHlL1UzikrA+AROa8EYrkchdhV7ME4q25AoK
1RqZXLNyN/C2DnMwcnfX7cm8wddFS7//2BzPL+7e90v+9Dd362wYwTqLs83qj65C2+abQEmTmhZq
4Dxe3LcxHi/L4Sa6VAd7UfvPLsB2NoB1SIPEoCt1EbLJfGEVq5kUvDRa1OltLqejwofzJ2CbxqYz
LddRUCLIMbaA7W4x4Gt8CpBt/RI2ThYOVIfiF+kh9xfsno1ghV4N75OFHxydLqQFjxdPxPkHX/dD
vIw5lSqvnTIpI1U23P5BV3fTpU78rqYRnUO9jACNQMDniywf0FjTeSfaWcT+phR3Ck47ufovom70
qj209/9GvC6P5r4GBq2qj1vP9r3+btIhvPbnUPx90oh8Zg4Sp6TWV9SFcuNGfP5zNV/Va6+YaPJl
YKmUSpVJeNUbXf03aKLxVuscFO3DXN4Z+YEw2HFpMZjDqfN4+U3/DDhtT2hI6M3swJV1Ut+i42p3
zI7qp6dIHI8O9wNqWsqHKHX4h5BuC7PXEyiPRpyrPCQdbOdKBV1Ku/rIunKldxEoi9vdc0DTsTc3
kvpwXhAKNffZOtKrxGDn2EexF+xE+gw2/WLXZCJ6H0KNtxOGJuMJ7xnX8HwPmg+TAUu11zYi1ZVJ
+ZR2dGybe048SwBJtRRlEuqh7Bohjvb02SRHi5YFsLPEzXGaZ/N+TC7n2H8IMLWR0hythZDPsdw+
j6KhfiSVMIUSfeq5VrOkCf/UJHHG/urzUpTDXFI1s4ai2BXafpRqEgJf/3U8BY5u8uYgg1etiLv3
36uD+/uVWf6lCAGBvT18es1id0RjPRuGHoyYdVo/0AqK6TLXtjZ5Da+yzgEPuTfRnOevgp8Fc55g
7afn8zijDRCLnPrc2lyjB0k+hSFKzwIS6k8gaNbmfKaU5gTqVQXjVOSEtt5H+ECFfmEARqybOht9
U7/UKKzL7UfreJ6RWmbbUK+L8QHEAzsIj874MyLSoQGY0Y5bX7IRvIe/l1BnM0sUUieqD8YMaKVb
hudFdMC9t2+G1fDD+N/gG9SlMaBO9XniplffF/DvC+Igo4ApscX+EkkDUCEc5Zo3cxGnNxOyvtyp
//XFt5B1ky8ZouxqkCggNE6RYdJcbsSkuOwFfLOdGo9vcAr8X67ChHRVhX57VtphWN8kg1HUtpBi
4sJBkFJmEsGjPataFOGnyNtPt30iNgihYNCCJTVFATrKDYSjtlIR1q6huqNBvGwzuJ9ls3F3gaJG
YkHgSSlwd5I8+F/cNNjANn5VOjGMeXCZBFpjccnqifOLhXUDkuvuA285gLCG0McneCIBsLoARDmG
bXGTJ7BlKJLIyym131uGAMe83/Ch0nmAVPUoLxgX+FMxhCE0FCy5xQsKF9dHxxcsdG8oHfrV4A45
8swXmvU5e6Gy9WKKF9eOzCIXdzCbYow9xum+ma6p6jk33D4W2/07/NrDEr6zTrjV2z+Vxh5S6Ci5
hSLypwHsS2Oj7XwDYaSRcut76YB277PCnO0Vez3D95oe1vsYy5gdGfdbXa7WpVuH+8tiTEiBVOwX
+/4X8DjmxjWr0sEYnBTux3dDN3feOjLadOz/A6L7GGw+2zkjl46XpMRw+/eqEZNC8qt7FOHkDFu5
b3gwOgpRAx7G+Km3jVNjtFfCyFZjci3WY2TdIzciFlETWy59KzOT7A8ao7shrw/XTsV6DeUy9E9j
48UtBUnSlpFuHs6uoZv/3GAcRq0aj+82s4P3l3kyjXuRA5kHBz+/RVN5/VLeVUznQUA5wjs8rVpW
Ti5z0C4+p3JRpG0wtmgpmCxit6P60CRFCjDxq9bqkqNGLHMQoPQH2Irj3jOUmUMy86vj4hbork7J
8hShf18XYmK8egkrFc6TXmMvTcQtRnlsCgJ72zD6H12XWEUz82NZKBfLstFxbm8KHjUshGKxe0gy
9e0cRNdbXqCV4YOZ02viz+8DPqLktyraZYCgamlsTBQxkuMy2wHik7oxXC1DRWF4MjyHyc6aLpFg
b0LHs9Po9P1ohu4jFSVCKsuT72EJ6Vui0lMW2XKcCnwhTttohKaYanXAdZtjpJsmJbpyIQvvJcDD
sMdkzZACHza0znwml/73DqYpId+wSvfe8QLqVRVtopwMydarmGgs5zR64emNwggM5/YAg4o+qcRd
EEzIyjBL31q5eR1G0EdxDfv5DIfIDmTPcH/fDpLj9I1hSS7HY78zpmh3J+r9ymXXfupES2ZQlool
a65Ykn2V3ztKJulQCOqHgG5iie29Bfvk0cxcysnRaN6FMicS/R9SHTYlrd5RIemlHm/yWtzg7y6L
oFhqAquf4+onrXwHKuU8xG74CYjAg1qkwzyaPt0jql0hjsRRzP2ZL0AHEzQn0OfXo4Cs5XlGvoxR
UaVPuHiIiVF7AgHFf7xu4RGcdA3TNjx6FMCBUyS59ysvNKu4KIjQghB4q4OKGrvdxZ8GFRn4lp1v
+Jd50N5JyfHzYkwmb7IP7kRwgZiWXFsBJM7czWfQZvIe7eQdu8rbC2md7oRZWPvndxGMcPttFNLj
c3MTaADdDMyrOSykRBNPndjjUfY+r5BpsCt2tvNUvwY9HPmJjw6/0clNxF3iJM41jFbEZwvX7BYD
8gbycEa/nF1zwpTpxkl6UGzsAxPc64hSv7mvQBDw71a48weUmNABl2tRT/+NfpxQ7/KJQ0Vj8mc3
BlxVxjaDMsPWWovcZWQqFE9DVDbzPey1NJdLLxKAFWLWjMLsyHohUvWbDPPCgvtepde35MNF8MM9
dCa/5wLfvpngCkhQF15If3OdMTC40cYuU28pX3huLnos11St6ss7CWlY+dJ0lHlrtuPxsQ1KU6b5
E3yZxO2yVqLOw93VeTW0CrgKNOabsaBjaNAicECOhJMSpln5NsBU+EAIWpWyXfuanbLnBp0KP1ON
7qjn0ARisbqR7wY3A2FUfwoJCCpfBsEAncFQXGavavmN9XSgRuZFOKoipq+xPf7jqghA/CBRkohM
C2tCOa4PnBexFx2Lzux7bM0s/UZwXwdcOhqvefao+O8jratvi0r1CR1R6KHDcBw7umed026TWfSS
J9DuzqpIwtzi4gTHTddPD6vKlVkzZhGH2c/ELkGE8vubtet7FqKMQ0gdj4IP3cGFQ/F06o11YwFK
iePFxS0qReJAc0czoyUaY2aJjpv37ElI9/mmFj6F6R7ndcPxlej3pKSomRRLxK76HHUeJH30fyMN
evNUJlD6/fRvZoDQqIrHYye4UHpkUEQORg7LferK1e37W79fr+FpDAgu1gFtiSbgG/PqoFNGAr2I
/AtFlV4aRvTISKTVAonkE+QPzY42EgtLesuzfXkhatbUcAXb3cxVCoDN5tsYmuaNxhAJdqkLofbe
T4XQdktP53VY53kALoxGW+uZeMgAExl1VZijCTuJRDyyep09xI98eYk6a/kiZiGuzwunVQTScfc2
pSWjJ6cjlO+bsdBHCI7Tna2jlKdc+lQjZvwINgC9iIPaSrCA/PbkPNbvjW+tpc5zh57KGBGlxFyW
odQ6CtSW/Nj4YlZzqyh1XweBwgGgYIpoM/zH5yiEFNSFr+TtN1JUov9Ge5GfUIpJO9RbqtmDmVsd
NZrQGzHaz+mJv/irLyphaQ7MFx3GIf2sTob2HqQ8tnCBVqXA5gl+YO8pvXF5tcxZJ7o0nANioyWs
7V7pUbElwXtUcRQ34gHFQQsLbCach78pVtP4yjkx+KP4iqGWIwbYRHVbo8n/cfEmBifGoWa0iShp
KeorNd1z92nnGki5xs+IWao0e/zWpsc+61SDbyItMX9VCiKCO19Dt8dLrmOuGEKtVe3e9j/40qp/
J+dT8NXUwyG8rLk9iaHoBRXdwQvfNai7BpTdR4qylJG08/6vs6pKP/hQ+R7g2afZAieBFnHXrTYF
eIdHQFs7ZqdthqDSkSEvokHjfVxk9YRkfWvc+mdznvJxlLFAFnNdP/Ww7XPzXPBqlraWbePNtsr7
5FAVGAKDDpcwD15Pl0MtOKhdER3De+EA10yT5xjagn31kzLuhawgRbRQzYYAB9LBbYrlRs3J9w3P
2QEYM5OsoHPBA+aYGvKMKTvLn2DyYY2l/bXEyTY4jOv0ZnP3sPJedV4QhuqKsZq/9oXigw8Kj6MX
vJH8Q6O1wJ0LRgzbacbGx3GfM4l45lvugTOwimlm3ny73RkGicvM+Bk2+Op0yLeiD/iRyL2Aat0/
8/9uuOqYWIgRbGq+rGl7mMaQNjZ3j+zOIlXq1fAsVYrNbqLMxvilSjOmGtpGPzn/NjGe1oCoxRXQ
AJgaMfXqVbfnCFdwfRi4ZgCLMzqRzGE2A9rL+oRnRtrixog8ez/wmQvd9v3NR9DE+fNC0kSFNAwV
z43bnwQvcX89gVPo3tM8gKc1kpCNvcDYMnu8+zxwAScjj+6jUh7IIlI8XF6zD0hKcu2i9DeQgmEI
Zym2CT6J+dJCxqDc0UM845K7V4r4weeA85EjuHPXXzLWo6Uww1xtIjlAPxUK0YoFINy8QLFH3pp9
wX6KsEzq+EAxn2m63YFMJfClu2ENdIigiPANCJFWE5+w+aoMhThhrW85WU5YjC1eiOGONaI7IWbm
zIPiQ7Lk88xxaWwBHlpMmSB34EKEvme123PW5m6fO56P1Yg6Gd+SohdGlV2nBGSsvNJyaqBYLZ38
CwhV/eRAGF+Bfk/F+arR0kGYZc837+iFvXOtPXu103Fa+vFcwFC/PpR1oF6cjpu5Uq8g9kxZqeox
deVTM3WEAn6eeox59VdLR/Go43q09qBJZY4bD+V3gphLibns61LYGSle/3JsM84Gwz3fM89NmS4W
PCb/ZhZMcE2FkoDlxf6dnFgF9HVxnR9yJt5YV4sEIS32R8kYgrPAF0xCZdXMM108IH+LDzysJC9n
kCbUvhPBUm+bwZxWdZsaEUtw/7+SUAESbkt/8V1paF1QRWXCMYQTklZgYILq9Urp08C7EBiTFavf
rSvevckBH9EuX8kju+aV9Bck3QLgmBMEkLaQqn4VIFLifZ4Qw2kkMqLQ08aFL5YhCn6R99mi2zf7
R7DJQlJ7KaZMoaRhg8tF6KG3QHhw07Bi34rI8xXaTr4PT5qUMUstBoZY46CbNFP2If5ziF3hxcmF
GAW4s3t6yZ46tRtJ5UouiaH6n+YEGHA70Z/armxf/YRAPds3WjuZ4gKoZaD3NE8bRjOpRcVhH4S1
4u7StBkxP62xZR3DrjkEyh3e1MqpCUgHgAHTG71C9RW1LZ0r9t8JgxDW5wA53+UmQJZM717uY7SY
S36ua51m4aj319bKtCyyjM+n0vHrDqgtEQyTKE8tglnvbhQn6NhuWtlJwmUwFyu0Bjj9CPB5sDBu
MHtbs/a9bWJQa49Km7n2gLZBU14SUVbo7VIuQbRCDHEJlqBqWyveivR+AP25+t/KDblbue4J6xnk
EV+EEGne7pOiWlRVYnGx/arBD03cL5OFcDH8D3rA7qXuTiKAWvEciMTvvhokx2izqI0FUUp0fcF2
KYL76JgXnlN9sKhkUMLD/+B6jh+INGqo+uQ/am5hhhjL1Mc5VRq+rTIWKiznPcDhGUG+yf8wTQdL
NQNqaIoh5Sf23yz7FpMi/Ky+EHIrwg8JkEiVTX2LKr3JKYGavHVGAGRpBvApWK9izM0UhwHSnmdX
lE8s5bxk1lFM3Kaq+8MsU1JpdR3u7H/WeUJtsYPC2okPPMqv6iUF1vt2RDxzVV7R0PwNA2T1qTG7
ItgTKZkbC7WOnkarSxKqCmWfFFGt7R3b1RadYkO0wQzGDUeqE7S0A6SUeDyfhS8ZRjlZvZz/zUPR
LYwR9/Ivx58FmGBh91Cbp25rh3rnjRIsLSYG883CzbxtAJMHWQocAwDxM7blPOBBKGYzWU/r8qIe
qSLJfpH0qYdlvMWihAD4pLZ0OASGoZxHA3XUc1O2fWDWfZNKueJTMQpryhVwfB/zyFbEtPUGg7hJ
N+5Qw4aYpx1MYdVqqC8gNuS1ojFD8wb2qsIkJLRngifrWMVlhnW5tgwMV/Nl8W+//8dzS7f4zJ60
V1VJgVmZGUr2NCGlG2AZ6cSbeLwW5Me7wLh33u4forRIcfT2VSmkRcp1gwfsPtSfdmbLEm06GOAi
nbCviNyUA0ZYBAO+LcVdCmcU3BOrLiCU7sQecuCJr3eKpZweUMoNWbJx7KBZoN7o88VHQTlKf+j1
ci0TPSR6iwhe3Qun49m+cze6T+wnqG01bgtgbmxH8dBLepLWwgNhM9GHePjCVVqu1Wz+bdY8Dv0y
i+LhKGiGeJLPM2cpFlNC1At9R7IzE7Tivflb8fLIyMyRl+wvPqzvzB6PUF5MV7ScCloHVf79wvFn
oMPM9DP5fXDjFIReVMIEIyoGNTaRawYy4hsTn71yjjHCDcsH3yKpW5UYmHk1qPznch24d2JtreNv
wgNpaaDzZWtdm1xCykAUHh5UPkdeZLCSWfF9SItN8QY7yd6JFZKl6E053TqfhSJIu6yWvvkTc+tx
DHrjss1xzWA4yOUPcQcdprhKHRbG87WcQnB1oVvvvQxO4ZyPtm1psl1rPeizLPjWgSXEsS3MpnAV
fBLpC60f2FnQoAnAhubZZaTAHkjCirNcgA4VuWlLliPRWDKQbpn75HNYFC2pS2rhLLw6jM0bZuV5
tifunjgkc3HcyfYOuYV/sHageQdwkxUzWqwF82RBlkm2S5ZBVePo4Ahsw2ZaJU9Mi3xjud32pBJD
TWX2Ngur0JwPQHgVrxp5Sn1tDgKI0qsNTKUaMnH1wn/u7nz6PWQuay9jvozY8ZAmH7prqcrd4DMN
h7EfYixEgZQqqMq+Ah+CHRyHsKIifv3cjvoaJGcMOUrMesmRAR1D3N+QBJG+21bP9CRv63TLfXkw
hwL99pP94lNoc2zpRl94piNUXmsuAD3A7T+E2zM+KOUXIaG3gjvKGG3CVZRvxmCH31pRPymSJzwD
9Egj9M/QgTliHAisNq1zZ4P9awoc2n49zGgZy43IcsVSr1YD/xgYOEphK6fOmVv48mr35yBJXOtX
YMjZjdWwph/clBvQq8HSlvZQimZxT1HOYXDhhfU/gTAiHk5L3a26RuIK4FAqDu10wH1U3scoZpme
rVgSlObfz6eJZpGYa0hlfnQaIe7Er7cpUbjkNIxKhPLTBHe+vrnNgo/QLDfyJwkltAu0v6uVS8/5
GeTV7Q+CxPJh28trrEoklvC6BMmVkMCPHFuieFmTrys23uFSZL7YRs3fTKhxvefWnlXpfxszjTop
ifYP00Dy/yp3G6xFYfx/JXov0y4hxxyrR1Fuh7+iE6RHNnRtXkbXkuz0pEyq+k8WypM8IvbZjKRZ
FRh7yNHuNXa+QoVbO+xRxE8+fVDtB727lqcpLExYD8ItPE23ETq3NWf0QnejVRdfiBjdrslMb1tv
8a4nzzz/AN6uhLo3KrOmQFEJpSCTZSBHkB0gjv7sqzykDvzLSErnoilp3zp5QsxqXRrvrlEBThfR
pdaPjxHejxLyGJPVzZuJfI+VfNBVE+QAnnpSMwNji7LK17PtD2z4vau+oJ16JH53fAE4fyjEQS8u
CJZ3LCIuXFJ1iudMXihvTtC+PO7rjAaPt5qcv7pWPVFzIWiI0pnOQukJAp0ItoySDINcDNxNjxaz
C7UgOecOpRJcCkpqfaOyTU9neKtec17VJ7Xerof6Wgy7VVF1kgT78SEpifWqSQlRxsF3u+biyUG8
7Y+7KhM1UpHePiHus/AtS89Up2A2Ja6y1eRSGe9fKcfXvqEZzKhXeq/gygqDl9heJ6+plkke1XyX
BJMapJ+fVUOFuRSGnueMY7901DLqGpQtLIhtg/drBMFahWqSM9UXhoca0zTkLwcGCUlDh2Qsb7qk
yHMO0lGgjwPPohTAZArz7nvCFRaKs7nhtHvHYd1zxdi4TqZu8k20287Eg0VIZbTvPuJPDCooyY76
GBLxrrbMahN4Jb1Rf7IGkwGNE87lMDxkJ09/uWMWM6lEUirJT3OMDaJxKNlcm+axObcPdauDghFD
H69kDwvNLBFLQWFZIHewGlivBK25mZ6KDHY5B7OCAz+Je0lNNQG+khLh3+Nh9xaz4q7D1NMW8Xay
yWb5NWxq9DrfUTUO3jtBCTrGv0AOE/MhOV7P8ipDpJdLF4ZmoAYiupkSSxFB7DBxMC4T9d/uPYth
HWf6DeKC6Ec3PXNrujkV+3juYAh44s69DkfPiVZ7UEkGls6hWpMtCK2USg1OzXIRvtLz45h1vBau
E6w8JdasfKe3zKE0jH1fot4mgIsxKzudWhRZiWnDIHOH7RpLbIUFjXhiKbo5hmpjWHEmxdcEXFSd
4uwHVnRiHvz8QbpD5vbtdQK0SAY7dUfPWZafjq7w8Ygy1aZDX5sZ9xzLLq7RhqJag3dbW4FIZg9T
ldb/mDfC0p2f09ueybDg3/RMc8vRQ5cmvUyz8mSR/QJkyvxHGQlEslZ1CTnA7+myJagaeDgjETiJ
ZOtAywKUVRUbL0BjLeXudqOcrjlHk+pS+cKLWHHAbCr6yeqNwMUaLj+nsnp8oND4cn/VKWgwRMsV
1VM9VnE4jeUX5/rUKapAzbWSHp18RRouEyKOAqqvmTwkkU2dYGCiS2yiTjWZuN6LpA9YwFv1uvyQ
E4VHf5NwVpA5YUDgspXQt+fb0bfMEizIVrl7mgNlEkRqtz1LHEfgWt7DJBVzIu7JxUt2cOTTe3hu
Rm6Ir666NCdN0GG8s0JRgxtok5V9TAdPeBNfBnuHkv62Z/M89a9KYFPYT4QSisUyaQUrFU/Z+QEG
tA7yZKgKEQX5/FkWq7iVvwTUc0U/4H+wSs2kFWUIGy8uIaKzRR00KgcyJjZbUk0lxOtaRbne3YXX
skijFuW8tuE76YA1gcAfvIzaoFWZIgS3oqOjZ3glCVVIZ3/CNLcfzhqxj/3sOxWsgZX+9bbBwYvA
7SmdgYOefzHmrsH9K3EqPFNFhGxt2oidC1pAoZwewilld578S7zi6gk3gcB/DiTcP+JwdDLGes8y
gXkX6ck9sI9EXBRpOR+58yYx95repLw2ftZX85Zn3bKs1DOHa5ZtFUBLDqvtTKTdn2odxjXKgRYM
sLjHEqO2J6oE4b5RkFG/Ra3hUQ7rNpiKWZgfyZPkpBc8Z+GO7cGSsPUdYq3/gchP+82lH9g21Szi
nq1jeGprCBQLlZ5BXVe/UKqLQ+jDcpEwmU/8okoQjudRvNp1OQ30vcEW0SYXNMc+nxpktLzgiN+e
TswhpNh8t8t8je980Zm2j31yceTY7nQ518OZtXcO8yipOvUd7Ri9wu1ZzH7SS4UYybZnioVMi6ix
1G/cFsISRJh/KwYJMNafiuMY7j8xe0nQ5+gAvG7U0uMxktttGc6juYVFYA386xPOH+Ka/N12zYTr
Rs6iWCoOL1/7Pd7z8pJYhrmLPzGEJxtJdbDrb1N2FNCBThTUI8fuBa3SZ/YwZnxUHmup0AxwMCiY
qtlypTwZgGLdUWGHGuiMBLPVoHVBTT8ZR9uHe0BVSZEFG1ZzTRxDoRI32UoFeumNmkaVnOk4tGlk
Qf0MaT+s+eS6AiyLulGoz/oB3qOxjlE71eOuZDnI+S0piV3/3ZqIP6LiY29qypWqviJfmqv6ywXi
hfmUPCEdEYbsFRvf1ayI3vDhQZwHN1GsK8B5YBJPDSiP23lpY7e/ihRMAsxnXT70oR7mjRQgqXWU
5QQTcVLvKIYH7pvGOm5Im4UorpsCwJgCPwhpSNVaMklu/nzqUrZe+0kGh1a9jR9zU/0GIEdTFF2W
KWH81TgbqdnY0Y+DMaGZTKwDdEH+baksQz1N9SmnLbFeoAad0ozCqy+QDB5vkuOVrFz6KmMt+pAV
tQjyLHbOtfmAkuKvDVvCbfqorwZxKBY1y3+96Pe1OLv6G9jzpHR4nCZcXFUP7+sewJrCh7LWN7CJ
gk+h8asf2zTdRtSEuSlvRVkd3kffGxTTeDwCYnjPDlyXy8UD+BEeaWMri0u7dgIIRKtQ0QMYV2Xa
u2exszhhkE8f1P4pfwJEfMAJZMi5VcFLmMX1dsqr8UPW/O2pr41uVJI8JJMnmo+yljTOGfRFQ9W2
gfpj1DWZBsi8F1GO4mVgyGlbL7pUk4ph0U9+FtfOfnVMbEU5LsH3T6KVXrcE1sEJ3/acLvN4VJop
/aZaonjrsfMMQH1sHDdq5AX475ZNhT8cRQ+qAWDma/McnUp7Jj36XXsE1TXTcne+yDjKMyhfmZPG
Bz9Ia2tsJgY8LFS1W0rzD1SlDTKKG3Xkk7bWl9HQzb4E3TIlFgM43++6Exn6m2Z/IfjFtCaKiDWj
Ib+tcgL2oJ3/umQ/hFmXslu3DRo+7+/63rT+2WSyDnkv6247d0obgvi/ck9ZAsXnKwwx9K7Pqa4l
OcxfQXW5AJM4+rdm8/dMDJ1UWysk25UmxUAw+zX27s0urMKBR0zj53YhVFMvvaE5Cqjd4N6VnBnD
YvAZx/Nk5gCYONf7TxfSSvFZOdUJzq1jVPs8iwPd6nJJHlvkXD5g7kNI8sFkhceyhTYaJkJbRr9r
5gm6o9hXm32XVmip05Y4CSErMY+55pQkkSrqXREDpyAY/+gYr/N6zh6VUVIdRZXJq0DsRmgaQr4a
ECXcH129SSDyR4bLuSePpRLAjBavnAeO3D8RjZIvZ6IMQmaFkYD7t0cJXUp3IXEkFGCc7eq0pATZ
luCiY98MYftvBlWpcgP1MVpufoYAAdzoQMgXsIEfYd+qGwU6NS6Bcl52GEh8xSAxmrdjcBb90UAF
vcL/UN/Lal7S4LDSkK2IFPv8bY2nzDzzh+fzDhXeym2yDO+b40nq3Xy0WeAhNeqCzN2QpH1/2qJ3
+CVa/WC1cOBa0Yof50dOuZoP534fjpzaKibOJ7mUHdoK7zr1fNH9+3S4gjDr4bZQKqc98k8Zd82j
Kr3tDGnCsJqUFiIsvNHPNu8XjiqIKr9UUsQfO3Yl8FvHy2XQMEdqlDJ3sGIz8f/4Evc+JrDMuq4u
jeI9XcvOLXtAX7bEdYfUUS30SRF6iXxXOanjKbg4ueZIRcjz5uUCEJrJGK9Ym2ljQHxk/zhU0ZAs
iTGoF7XxQc1sN1VWGYf/GnxcHhWGNROP1kOCvzxskvyuOKDCu6e+6gToqIM8k9VAv/3zuoeikH5p
Exej/jlTpBoP6zKlfnju3ptYjOBgISJUPC+uAa+vQRghK+mFcsjx0qMq9t64PvYuGurrOpOIY9fE
ut4B5yfHYVSBCQaJ5zfHYDuhopHlpYv5eGxRqYMje73pvFwF3yiU6rxCETdQjjFyw9SI8ogZTDbN
hnBw+wNintME2STSNDEQolN21d8Q/LfZfnYAo4jLQV1Ykx7/l+69jiPAQBj++Aq39Ju0LsmRMFT5
9uSWCCoKsJ+3H7gSAIILkqC+21az2XpI5n7KUwZI4m5Q1AMfEaYdL9w8BG4K1ku+OLpp1bTqLTJm
JxIzwlx02mmCub3VSpXY6yu3kWUsbdQyXlxon9mDUIppb9Hhe1zrWxckGI7Xl3pHPEFkhOSZao8q
kZIn03Vdy6njBQRi8+9s40iHllxvxQsA6IdkHGzpSjT+BSjhBPY0Ph8VLa5WLr3quBq5iQgtxOOM
rJPpsVd/b1YAauJ18Aa4fkVa2jLuqz6+M/orH1cdEvEolcqJnkxiY0+TGSbO9WPUwsnxJPr+nzjo
C3Wprn1dBgv1DfOI/GNRMm/C5sLZ/6/uIFFQefmnxna8EXWFYgPvjh3m187yNt7r3sBLXkaSQdyh
20EXpooaFRTbOfWu5abfY1Y/utMy0bH6eBxjwRaqW0VZxoKSb/5mXb7iLWoXCNa/+1klFutu5P7F
ROj7M3SOxd6PxzQOPkHVCAaYIU44OuVd55vIUy+7hLqozMCKBMI4zvrXnHS+YiobEJ1q7pIPc3La
QnIdCQLNLN8IP8fPFwfWdzfbMQMHhkscySb7/27VEd+ihzwseBvpTmSOzm5ElFjx56UgC9qAllxU
Hpj8OMa+/y5gczxlFkdtWshfrtJywj8yYnm2cAjNZwgdhc5yQfxyG2PGoR39I0ujohXlM+cJqawu
SDrVXiQbYYr7n0H3qEEctvfVZ/JvPmzWkc41TjFltEUQJDAi+a1YHgRrxdwGGFVwRfUbsaHz3u6Z
mYwSZLCXD8iy2/M2pm15Ub0adhjoGkIOGEM+AS3c+jF05YdKsL6RGZDoAmrVL1xioeWrifcR15Lo
bnsyDUvfF+okqAIoVoVHZ1OdrCfgX8d3R4V5IhscbOa240gjkscf0GmtCB96Q4b46ZeJcMUp4iPG
O1j8NaFXJ0LHS0fo/YLHFSC3Rgj3jq6GT16dHUMYwoZ2fcqRPC2F7p3DcqDj6cBjOBZqMhsE408z
/tbZLYRCwqyM5tLVUdqxtmwK58r7srZObxWhF80V6QhrUFyfb3N592bBdz03U1sENj78GDRw3nN2
VtLONq/rMD4+1APtpKG6RPjKKK7ysU8vaKMGoZcnm0M9S86Gw5jBlS84WShdIk6xg/6GxM4pJymS
Mb+Ap43yXmGEZLIDjrkolNfXvz537o2g9w/O0+BoX+qyUa+BkquaA/zkYbcgB8nknSQqaD4htRB4
nt+pTsvLc0tOZCRZb5CHzSHRYX8JK5IalgRt2AEMze+zgCvdedGZGlbFnJdgJeGdzAggECyEpuZ6
46PZR0ghhi5beRbQ7+dZpntgLg/RxhhzTv9s3MOA3oVPG72JfC8AZSijGSDRvR/rTY7+thIRJ0w8
k44gFjQo0XGb+5yV/mOOd6CGDryBw94BfUJmy+3I4wC1b5xuQ2+8eySpMr5rNlAsWSb1S/IIBD5S
E34c7oXwX7lyfP/J4Zj2unczZCY0FddcIHY5QH2cU0tuT9rsCqNgLm0kixZGvGkEtCw+5s/8jhwE
/qpf2EEZVlXPs6ygAYVj2zPFe7vTgtq6WN1WmaxktTxT/dpZr/DYI3+CT3bct0WXfhkROfJlquX1
gzk0E9AdQ2EUUFKDOcQJQGK1kCg/BSW0e9iNwIXEQ+aE2zJVc5T0iXVq9DDH99/LuDihwimGpte5
zbPKPiVOoKqhTlqFzVXZGUczpampYB8Xc4AqFWOXX7TgS6w+SZUC0aeu14aOUqN9l3m202iIwuBK
WBYnz9r1/b/0peszi7AyJATjNbDsT4Z4KbjUKWUw4lONMEw9CdswLW5JRfcn2UM4a5xT3V9L1uok
PXmQbmCSRpLMD6XzszhU2IcltptcYIUa3v/MZ/YcqC1HRCIYOrz2ERq+s6A/0yVOGO2WCV99sKc9
sFxet2U5bCz+NpB3aCz5ne1wqwDNFk/h5nXNesBN9uakf6QZbgRfxa/6CA+iuo/JtySa+kCyuJgL
pQH1968CSgRy+qpgLR14IaRotpvvy/58pWfxLVqA4eAmXjwY2ha4Zr+xgz3nnrn53hy5MOm0GE4w
aVsnN5hEKGVvob39kH3e5+kMLh6EA1rhkysqmuwR6xJ/iPRwlBGGu/zp/l7d6GSULlPZbWff88BF
QOpmJoATFy8Igrci+93KuhjEeOGzTlZ8u40/z31XLAPY3OaU78M4aCOGOWbnGX4J7o5hhc8yOqB8
XqRAw2QxdsCib9iMcHHGzrS0B+L1QHf/nkqqGGDpk4gJNOMUhfcs7KBjCfm8ZxEb9sJwwyLQH1Oq
aXk25uejwUznZ9fShqIK6lj76BGQfyWCbYQNW6hVKhf1NUBXUU2tsRx9/SCQnC8YqOA6FOTdgm6u
PhF+9sQMDARRbekG9sj0rYjgsfZLrjJu7UG+C74GKE1rilGGyPRuuBn73CwZ19fHFHowMZVYHDIv
kgh5weIBbu30JP6xQRC2HUvyat8XIGjkI4GlV0R/88lZrILlcM64PS2mrD3SHsW//xbx31Bz9jmW
Spk9QiHA/L1xLQX60h0CVQbMPkssNjZgnsL2CiiCOF0hI3q3Q1L5eLCX0sO0ImOa3WG1JWVopfg2
jA3Kv/PJaR8q8oXm/Tu9oczDOBiUj5pbQ5HrRPxc3v7pbC1h+KAS/HT6Kmz87qGO93TBZxDW4PpE
+nkUc7yvnMRXMJGCkNkKkGyaXtlRR9SzeHXp2oyZpAc7OBM9TFgAm5kLpmc4iGxA5TBGs2R8j0zp
Q5SkbymIPhJDTOsW9PIHSwJxBlrJi9EDlDtSg2P1ZD3pq3py0uc51hJF60VnHKCD++MtRS38uTFY
c1V12Yi8Yqe7r9xkD0hYWO30sxKItnDw3VwsNxZtTSGFN/izlEoWsi0klCtoXhcw51fUYwbzcazt
nr2QoU16XQcOjZDMJe2rLm6lpgrrKha8GPDOOgGAWSU+2epN9fYeciiSMYd5HZHQLt1JXsLlcEZ0
zzgyVFNkfqDRBCqpl6r1hdBAglAanciIY5pWEuG53XoOQCf/YNX4a0TSO77pgyFafCOEtQ9MHzul
KBi1H06ptCNF7yUcFhDKmLgxoTVN235xWYPEPuJEN0/3L1Wk2iwhtUbQer2/PFgxYaZtKc1xw/fv
DhMosssB+lE4B19MZ73iroyEXGWN29SKVc37rtC7DwwoSPuDPHMj69Mg86NHVSGFjqszp8CLiQTj
Z/1BlfO1nUkNdkpggE3FG8UUKp/C69UeVh/uhVAles2C0ff8igFexCVZeZ20oKC+kNKupNne9x4r
EKhkQhdKyYphbwd0U8H06iX+mwXsAsv2C4taIyulRNRqcPj7StLvVBKEhZKLjrPknsrdomnbtxoV
BJhmgpC00k06sedxiu/t5nWPR+l4OvZVgaMq7JSHs4+QFnw7mXQAVE4lpWjkZaIyFuI0qnle9qGs
UQ5BS0/asp3Yzrz0MyEJnPMrchQP1dA+VQgGqRlJIseX8GTqw/wMD8Py8I+6bgEvlafIDWNaU++1
V7tT7Ghg1p1eCXGFD13/Bgy+JB6aL6BC7RFQCRR22pAbqjsYSDQc3tP9p9y6oncFZkh6SMo1bCVd
103v9eN7ElyqqMl63Jyng3hgKgAgK7A0bBR04W5Ta8S+ey0AbP3HFwJ/WzGFrOBds8C7wU5H9Ejr
8NDz/1esPrMKITQ1j20LuuPN6XDEJgTAi38S3kAVWYowOkRSXeAbc24kLJsixdwKcNHcQ2GpGpw0
R1CyUA+Ud8TLdqsJwsHVpgdh5tcuCumQ0pCoqoT6pMj/W733Juf8jWml5AjUQ2GGbT9p3a9cM9lw
4muzs0cfdxwRc27MlkzERBrVtYP2NnpEj5RtG+Kaqky3XN5ufDjzromjvRH7ECO1O4INflLnuaRH
MLCjNSoa/YQBj0BcfgZG1OE686pAKOjlHuiWiFJ36XxUV9ztdNQqNGTq4we3hxMfqbw8GtdCmnFL
E163uQ9pQ2bsudoCA832rYI+w9ZPvw+IiCcrcBu4ltxGcC/Ul+183/mVhfdyOcksb6saAOJJNd64
7BLEqANbsMGF2pjOSw0e1KvNfOQJ7vabB8s5gaHKGLbohMoAA+uQNdzgJOmecFIV/nR28RcAJlzj
1UwwW8rQiaekwDJ4bwfc/Myalu7EPrDfCtnCspKWEL5rFB0ui4AP/6bRCv8fhf08Ihmeci61TUjQ
3C1zONjCO6qJSH2edy/t3uzGOdxblJUqZ9bLZ8F82O1DZ2pGywJICcv3nyiuQ95K83AuzTEEFJdq
GNRbfuHgP5PiNiW1Hd49j5xh/fLVKdGTERlMBDdrM17Z34vFrDLyuvJLs69xubSSd4JuV6kBpnFV
Jcorr7DWSHuhoKwlhJDSF6j8PBg5i0fkecOfkCtQVLnJKbXFR5pXeJ5rhJVJxBzhvLPh2k0imOpD
kjRqxU9YbnMDj+EPCqmUMCL6VWfU3ktf1tg7v+VyYoJ4D0bt9N7Srab+LwYrJJEOtmN0Olc98z+z
5do35wTmEXQdiCE3l5OdPp8W8EEw2Lw9vVPSDOJBfkebr9+ZYxXJFHQmP9u+0uQomostG5yAiJrj
0Vf6ldJY2SgeA9eBglrDOFn0tzLeViPm+VYnF41NSNhB7wqQHe36mLMF7eqJ0GTg8cPvjCtNthcO
R8pgZhG8HKB0qNRLATIjGUmBx5LGRRFRXVzhAPTJHtjo0CQQrMy9beldRVkLWYNJzh5Z+DbqyJ6e
XvDVZNjpApurZiiuJVPwlSX+YK8BfmvWIiEdK7oJs1n/OtgNzJfFMLqDTWci5ZIokEdXN+lwSlqW
PO3tmIDOPhXVCZZHhToeB6bb28qO0fksE/ihhlpr2LPhNrx7dfI2zNu8iHJF4hqEG7xpXGyB8vC5
lVNEaVyT+7Y4WE7Lt0WUU5RsTfui1k2SLMYQsi6FWSqnGwAHj2VC3BV+J0vnkdxYXtcjMlwOtEgo
S9dBnFy0OHLf9utGOwRV985t2kmzxQp/lF5JockNGggtRtc6f1ePxUgzZa+OCO4LVbM0tal3w7VU
xrJ1QHzaXupf8zqyxK22IoEPYEyMkqSeppIv88J5CaiuLUmLG6kRTxe8Q+NvbcXLgqI83PCrNryH
Y/fAhfScVj0FYnBVGw0GxNeVH7yxREOB2rIRCDkl4UewyyehaRRqoqmBHpfFm3Jz3sW6s6N0+HJw
nMop7qd/9gx/EiioVm5dDb5baQHAz6OpaKqFVwMmETEC0EBj9u5OlTzfErhtkCvRIm2vTbmfFDkU
om8RVJgdryvWBVapNAHLrg21UNboR+ZnMOgG+1pWkBjhk/HNmlMwOcJNigSTmtGJa699W3VmlS3E
gS9nOUGarFxOt8kdjO+xOSVVIHQ4Y/hpxWJquVxgz9nOgmBPupxpcy30dlJHCX+r+H0iws56+SZC
kAK76+HEUxMhQyNu6V9uEgBarS/svDaSnC/+48esGhcp5HBZGankTfVPCpsv1DBtawBGGbbzeIvN
mp0+xwTz8lb5TNLZMB5Kynwl2Ilfc/yrOZktzO4VfapRp8CMt+ZTOXAA32cDW8NGSf0tbE5BCXN+
G5C5GE+NmaiLv0xalZWWhP1qYBPEJB5xMYENZrewpt4qp2Rq7nGdnQ87u4tjaA9bfqHpz/U8OhEH
y+j9Nif398MolnZ8IoAap9N51zoXTjvTkldb/9YKw4yy5yiq+qrZjszix2gHyFFJVpCRRPyYA5W8
SZ8qbxmOqBlV1bxTCPDfqGUSdSlTIxAhGgakNPJAWg08OHpyq2ABQGSkUmnJQ10tAZ/S8osd2/Cw
LwWDyvwXi1VzQwtukYprFj42rtBHMOrof019a0ZyutHarUHyR67UaapiFkzSRuetn6QWMyOthmcf
h72vIrUK0k+AX6llhSXnkLOYVGrLgIimy7aibhsNvTglCgstz9s4LcK6uVwoESYC2+VYuCOIyRfw
6AQEXxhB22V3/QFJg1AlpaF4ezsS1Mz8Onf3mA/O0w+Du+quWXh7/fuafTWzLQ1iblo8u5sWZ8nR
Zwk//m5BqXZPzw7aMib7uHcYsswTBnsaECSZeqf1pUx5uv6zRBNsSxh8NJ8xDBvhb7lSlaPXhxnE
PKmkEX+M2GogYJ7A03glL9HZcvu8tjNkTD2ek7hqWwKJVTym91gs48zA6RKUF9YdPITmKH+kUf0V
UVeIwSlFEOMHbbuICgHfPL9rCJJFBx8sm5u2mS0lQuPDuO7LekQXBNaLNKqnoP0kuUefll0UgXTM
l6CypglRUrwnpZJPBCPCaoN+DBhD2swCOEH8eC38C0tg/ULSmuHUuWgFuKKqNADNn977R4wbBty/
XUkH7LFke4uFrfXzWJAKmgoe35n73CCFVDuIXQ2j8Ncy6sUzhxscEkcLRkgnX3AoM+awZHnavCNs
o7r4M/5ZD1xdkUJFT+VYgIVwyGqQ6k31aOWc99IevADVxB9Zrxko4NiXdEWgeUfF7/w1CGENkuM8
EW9hA6Jb6ss8YyHgxZRMUhkoKfeKcNCi1xaaCJouQC7R250AmFJCW3TdmoFhc6GEiEyohCzLbiwA
3q0hZjIbXMybjXLmawGQt8ND+IzVrdZoWyHTeMWmLKMITZXwg7oK++U1ND9/lZQQWdB1g2pmkSss
SAaJ3t5OhDd37Tgwq4niCYTJHzYOduxjFd4To4ZVzMDKLQRWeDao/fg0qa7uZZ1BJGjDtMEIXKBv
sLJPaudIWDplimY4YEOlXdv/qYOtcDmybPyZnDXCwfv8BZx4Oo2QO0rrjxSXH8S9duyGriPoK+K3
X8xy+ZOrRTdn0lyKESe3o9i0B9irgRAzgbgZFcOvrejGvw8tNVyRD2nu28LdcAUEehZLfckUdef8
lVDAcuu3XMIB/FProOxhp+YnWXfj8/SVOL72eRTDMEvz05VBaU0CjPH1xOGY/Abj/ohci16HrHL6
Wx05yMCD9Co5CXajG6CD+/FxzC0uhMKvE9ODc9d+zWyK8jDhagMDE+g5eCI6eRT9N7SIDZ/91FyL
5zNHbuT/aVuRIVZuQRpZc+GHw7Joa823GdUa6B45GtGeuLReoG2BmFnY8VuI/qSAyLnuiVs0tm8s
Em8HU4zd6MGdwNj04EA1+62jY2yWV/ZVCeSVL0j2pozfjc9Rndq4V+S1q06t4jpTbT0JwwWpj0Ro
oOiyU8s5YomBRguJtr9R5AenVsb5nJ/KZswgW0e8w5VkijAMKyNbW1FqEjNkJH7obIk0v2NCrGPk
tr+orNPdHuTP5P616XJpZ4xOf9FdIvaSZ3tIBjffoboss2SL4apU+p/ZcUu074lhsw4JILJRbLbk
yYFcj75Vo4b8fyl3Rnp9ZaW3a/SkHZWsScfIO9B0XJfpbdZYQbYoWuG8VVVjkM93Ff/5kijt58nA
+PKsBywSOt7oju9Ku6MLz+Ek7k6V0W/JRJpvsA2INQYC1FI02i8pihsNzBPm/9K7l9iR4Fd0SDkA
wvxgRe1Jy1SpRlQaRYXmSACb3bzSr8HGpVz7rP5UMEGwDYdy7O6szmBL80YCpHJR4jHUODOjqVWh
gbuF2r5Fqqnky/eeJ1egeeC8xCvGmyLCnzXAHg7MEJROTIpwj6PFbBeMwa6y4JrYgE1RZOnOUKam
hkXDcQWZGSDgR2Zvh6UfNPuIw74VWZCFgjAmKY8ky+feQyXWyHZRKO647aAd7AndLJtGpOOro/Bz
Va9/HW/vq9jXR2m8SXFHnQJhA1C1BYBy0rPZjiJyH0Ts5Di41Qn7Zcj/naDbFTUvpD4cHb+EOgbE
oI1zUZpl68+8OB3muQbiUjMiPrb8XylLU67JZLKoLfkECdGImukq5pe7qKV1q5a0w3hZLaQZJkRN
6jJrcmQUylfUPcyh+36Uw+av0Dh1Ik8AO+8TPp/OX5m6wcs8CkYYBTH9HYSIxmRS1fQ8qJb9AQP8
XdQ+oqFFeLc3BKGyIrQvNNE9d5kmdVPt7+drINMwBa6u1oQwPHtT7E5HJW2RjJAN7GDLJ4AEYqYy
i+9onjZMceXREWZP05B5UqrbWos/Pc8UQWqO9dzttU2Qr8FixtFYEXHtQEDnVBKoK1I2DYo1RneM
JJgSF30LB8YNuHSVZPHCw/MvnpVy20Y+GBkKu3CcJPwwY6lNjovz7XxTEIWqrDSd1KoOcvhDe7yd
Hbjc7Xzqz8K0eDR//v/jRhWsfIw4ViCrAdhUVAFbeWEX2eZ3XtKFFK/U5vT4jXX0JiQG12aRiH7q
yCpBKkacPpxEmaEmbF+4MuVxpnjm6suGYvIli79BUKjEPLgL4HI92HszhcBXRG+9kJgeEqRdHp4o
6h1ceq9vaYKxdrEN5BTn6ig2UBmZXnxGF3LWqyPk2QQrzv4Xbp+xvFXAsa0IXH38exL4HdgbR7Ib
0pC+7JNFKyh/IC2atLPIX0JngxuCamYVkYOSVVq82qsa36q1SL3RNlEFEYkiWEYAlKSDdx5oIYmB
0BOcYLKfTCDLA/4hcOorkRkEAiHHPeEtvW7U3hd5GfNTjqAtx6vV3NzPLyLk2z4eAudqX1ZyzmGG
sDZAs4VhcqL9BUHKCLoCtnwA3Zst+TChBUa4GBLW0QYqVDY9frO/AoRsQZshPmzhPbM8moBrR953
rFYMX5WvZFC0j5XpVoX70UxhuVZdxe//1QfrifTSzL5DacKrrKqJADAAyvAFLn3q7RBPaSrmCKY6
LdKyyy3lwGztwxYKA6s9+mbXe560CD3VFdkp9JqoYS0RokaU3Fou3al2QnJJ79ECbAXrND6nwK0/
TvIVhHrPDC/Ym4CunZZlegPJ5JiOWr0TQ/j91RCS8JgU6BDWWeevq6qfX5Qouh0xbXJ7HpeoJNAT
ZR0dUy3gkp8M+vWXgVz2g9tjzdhyWmjcdi320dIM3xsXQOOk8eMaBoHX3ckISTiETglj/GNu0WFx
zkUZr0ukxObpedMn7lJISGfIkVE3dD6d2v6CIbJzEU7BioH9JH3KYLMhrQ9ycX5xChcCAI/qJdwg
CsWmQYT6XJXUm5IbOe9ZLvQCiVXcYVgA9Bs+ZcSixFQh3kZmSvL87hVQrOIYCYI/6exhb78N5J3t
Kp3WZP3dThRV88pnhPW8JXlHjUN5FpBxu9DgtsBn7AAhVFWgHGvRtIBeBNiHhP8O646AK24SabKV
p3jp2HHKEp1buybXqHBGP9drKMv35aAKEJpN4E8+HUslFz3SvpDojTs8ThK6js1IX21AZr8/rWpK
Y6D1KCqJBWLqbjBAwyEL3wxA2/exBhAHQ+wha73lnpkdNOzj262s/yDcX5ZIlMRQnBJk78XsWmw2
z3ICKdB4J25KTgxl9IEtcTKnC+tF/mXO5TuoNnTj4rADRIJwumsadzxti3cPnw4E8wGWGF4KNkt7
+BXJJi6p8HMFfkUzJlqVMKUiniuvWJ+BSNd5Y+hBZljAGAf9O/n8X3L6v3X9ydmdOetG0CsuZiLS
KGdvlaHHU9052mVktvj6cdaDxNjmNHw+i/Le43ooydikaw15myJB7lHjiU6LbnGTNJr2n9ZSmUhD
FXOxkJDluKKX/9oSXxdI22fTlszmf+awSaR8MnDDRkYOiJUXdL1ClOuBaYffLiPkykO9m4JApRSl
GZuHHpHJVqDjs+S9DohMT2H2Is7741U19V1tTDG63c18OK0IKfxinea0Eemdkc0gCQ1FEic8IWXc
7W6GxIMuskuFz7nE8z1roI4R7fC8QeivmEO/9fXhgr9gzPNhe18ThZ7sh/N1Gj4DqjFREP4EAW4b
RRcHQPOinE8BeEpeeGdv6Ar3CItaTrJ8SDUmlv/gViJ7WbIBkA7KGI739gNhv3TRW4dCGw1GKLGw
ceAmTFPU9eQZja0/uIQXzC472Tcekk3r+OvlpfkDtoVtDbkbT0mkbPYab+xOytZugm/mOVNYn+eA
ljEy3i2STK6EkV3FQFl07/sI+DLog+wegvgkcYzYVDIoxbB3I/nAStuo4AKbxNwPjM+NBIWbk4/z
k56AJmyIn8h04Y7HjYJ9sh88uMrgskdac2A/KEczoUNXrkWsEUrThnHK3YV55tqxE7rF9bGZMpqI
EFRPLDwt+Ya9WIvpZ6wGbYOYC9u1mJ57gJXIwABTofXhJjthUQXzMDTNs1me3EdKhL+nj20sE8Ob
tRMWqM+X1PueVgU1BkBi/f9ygxOystiNst1tIBZuScg2e3MLlFfb5/aTHhF9wSA9JJaVGTy2LX3F
iQQYgkgeCs6IhqYBziv4Vh1xpsEyUobjLFS3X7JnWVaIR0hkNuvQalX7kfuWHRmk+mmG/ydl7oy6
aqO/Y76MemhunGf0VQweS/eu/FD06czjiu35lGQtVNK3TYAY+8NWpVA2uQKCE+hwMWMlA+2iAD2h
24Tn2xD6cHtc2XE2yUtKPqftzLeryM50PQbZFXOPQSY5DSrfxxOam0u3SorwdA8QopGn9sTR8iu/
cJwUIeqKxCfPV2TVcSeUp6p3rMnNBruFp/96M9ItUnB/sxcM+6jnPh8bAzmVkaF/WInsGf99A8bL
uN4j8ykyypAEOqMvmYvguSxWe2rSkKt5YToVSH4cJmghzikEUsNSNqoVmH6W5aaI2H2xU+tvAUCv
HB3jAEvXjx9b3h/KYjFa3l7c3/zqbaET9Y6eB7td/ZrpYw20nM4FaJCML4CBXcZKvCUtIkiAApTO
6wuik8jLrrxdisqzJvGcTZRgAvSIfReewpkhC05FCOv5ZUis4UCFM0RF7w/O1QjHgPaaO9hk5nJM
8yP6qwPLlZQryWq0QO0QjCC8BFnhAf955bC7+i94kRDvgn/JzDOQXHNsBo+h5vr0AhlQgYvhEXd0
CvPTFabbMK2gZpR72YJFgpVLf0wij/E8NZIApBWoBnlhsIiF0glhZGXWKnhydrxYzufuxvmgCuGN
yW9t7TqtlLIK0gy46ROGU+raa5YEc/lbZUr2iOinJ7dycRRQqf1lY7GWdQMybLmu0a0OE8xtEOTh
eRfrCtVeRY7OP4KzNnC+hP9rIQ1cQpXqofK1nBAhsthdq1IRvxWrWbpL5DP7nI24WD5JJUMM6Npk
OHqpe+GLe5fyuW8GiBQTEgnHr6RZJ1b1nvfAZNhx6HnVoSyWcqCwAJ2UCrsN24zxkUVV6kO6sthN
XL+P8xRtsx0z638+OGWZG4VLsKCsGMRcyi4twagrzxZJlHt7B/Qirp21XPmoQnRkMSP8Sm1PEwTm
dSPBHd+L86usLKpnKIj2ouNTuLceliVlHFQInsoKCxWLgUsTWXOSwZS3nKwrrPC9fPM6lGAyo7/n
rOaothAqCvIRMW7m51Wd7/Yeb7uP4IubkEeI2Zh5VfVQCLKNolTeLkko51eqNc+aoOA9Ocs2VRrx
WQgyrVuclq4yb3umI/tn+rTwp2qCGDUTNk0GsO4nlt5EI8mUTCt0ncdDsY6HANR9unuC75MAIPKb
d8b9zwWesMqCI1VV3m3/saKMPoU7peSC0AUVyL/X51GuHEwZi4+YfWx1R10hKEdk3RmJ68J6a3d8
wNJLbutGE2b6qq9N/KqzSyH4EQLXJmp2dSqzqwDLXHjUtRj9JA9VZ5RUPN2YkuV0tBk3DZKFBVsV
AICDQ81hfaWnbiPZgghwiOBXpCtaYdBveOcktYAtaI3b6W23ctf59nJBCIsMRjK80N+YxyE7mUlh
K/rac+Sz6Pvtg1RBG518UHmylaO8ONqeh2vwHf0zjxRDEpIlW0rYO0geEhfDhxCl2Vwg5xExRiCf
i9+1k/SU1HWPyCgcloJ60PabG4WxTV7dyltwed+wH90fIBg8wOnRdYEPimRg6n/dvMczSPX3r1DJ
QguDZUtQ9+JsKOcCHD5vYiGWAEDY3fZkWMJEkNilXc7H0BCWKiMi2iq9OKWljAQxXORV2fxPnR+V
TorXOcnf4PCq9vmCSqIHVTvKZjmGdxcCxj84jgp0LBODNp4xXVHGULJut+R2aP487IUMm4oUmDyN
K/MEnYAtnz5o3Ydn7QK6nxUE75XDLU19FfBlLeIfAr1GFmukCx44NN4jqekFf8s1/63YwU/vBn+E
2L1QU2Y0pKtPE2xFnH/ws0nDvG6COJLV8qElgFhiV+xByjrhb+7wotHzGasShfoX+6vw6GcpfkXo
21JHQrvYb+i4dEPPMqKQmgVyQ5Po6dkU6h1pVLNqezn2fiXXUHkjCkWp8UBndLDjx+m+aU1I7qmX
tb/OphX6jhk9xjaoKwo6K8/4Hs1zBVD72CmXFM/j/GDJ3Qcl2uAa5pzpyOHT4czNmh+NOUkrymAM
NG2f881WpIWV30P7P6GAolQCEPQNfUL3yxXwTOpjoKU8gMkNksoOFEC5quveIAlkVLhr1LRjuTDg
iWfIGc8WaQAqsDDmBFVnmbR1LVXTb4fWMEopS2BDDxcdpuSH3KkgBuSQSRrzpm504KVQ1nhTkg5U
nfSKg5s6q5ZfNhcdz3nbnAag51nKtnwxIGURsWbNNjKySabop1E5uDMw8ZRfcxLuaEvGBPEBLavH
wvJ1NLjDqNIyaJlk2oyoxsz7Mtm44BumH4Zg8cmJOYvZqI1+SqTGjdf+TRtf11fUF/yZ41Fodztv
KQMSCX1BDV/5I5HWsOnP85Cp13eYlIo5MgSfTLl+FUESUGCAJODA8CfpW6hhvqk5I1tKIjqmzkm5
Bl1Ybzjnzw2JXKSQJB0/n0VO9I2PxoDZ2jvK9yf22mIazxFUoifSqqvYF75c3OqLA1dBW1cqU/7O
Gx6zPg/2kPeNWHdnhPQxkRa/EQYogZWXDJbjhtibxf9zuEiTKX+ivjMdlQ2ly65PJkzpZcvLwYFg
ABBsNfqJ7Q+wI4DzMfzfm/z4jSoe7+ntatW01ykABVxXdN0usM8YQMqzoG+CXN/oM40nD7BjRoTR
aelz1DFwne7sYcAbovYehkZbVRCjrvP2r6FPlDTHlRLM5ArTKOXF2l8GMV/Qmy7FhUbJvlzEFf56
gKNttkYhH2mN8/uaSVx+Vh9OlSJli5aovVYcWgcfIZ/5W7h6TG3YM9FHUoEAjeB0SrGil7VkXJ32
t6JudPxSq4c437XOaWkECEeaXtCVFKRHyZP996Lfj6cXUc/QpDzbThQxmI4SaTkwj7GIRU/My3XK
yBRdvLQlBGaRlh691g1pDdzGguw0WuBdhALxVvmrf1sG+oT9DfsG1/YRWgXgaPseUmt1LOiauyaN
NPxWdjK0vWibhtpaQFQoIegc1/WX5XLt+6jl5bOqweAt2g689lcpiKJIBnDXPid3Gdm6GV8l2Iu0
wDmSdb6KI60nn0gS0oo0XS9xRCCJfWwjGzLzIk2X2leAo+/hXWxyYqT2NHqtBdFvYhsY+OdshNHe
3gIMsS/BSjWX203Rxcc52qGk1X3WGAURmowxQw9BDbAlJuyH9pkANch7D79PUThgD7HaIyvBXUS1
BPEOmT2bXyp+OMJkzRS3tI2xz5PSHWDmfc0PENSOVJgyJOmW/qe3PsZS3k0pZntLBUuixndPC2BE
87RZJgMIufbdKN6/QhcoNeP/UcdsElD0VR2sw0FQPODkP/dF+ELqZ1ENHccUGgeVY3zd3JaSDYoo
4pDKDk+dBVDL1pB9i1m+QMbYVfxTQDNqWaFMghJR7EfR6JR1LwMUzo6HbvD8vx0jn9AUzKaqPpgU
gJpAuupAPio0u5r64EHjVuX5JU8K9hF/T9LNlLv9UKT5IknxemD7hIq8ovwzTyyxToxOzQqObIfp
k5DYI1BqdnrR3NreODh7crVzSPHNIWL9uUmgsjtJ2FpQ6qKg0ACQKJO6J1j8SZaq0hBJWN1mhxyV
d8S2rNjUtRMJKaCrtGCJNJGZ563sRoNk4PYDBdRGYznlSmd6qlsxoV5D0fdXRuGQEk0V9/Ug3Qgn
J9XxgFb6b1AwrsoqFKqqjnhydVC+FefS9RWTaEU9i/Vj+DZ3Lq9RwnJYwPavjxVuGoi2DBabTfd5
HLAaubfXwPxHjThNqxsnykCLEQry+hMv78b/EiDeCCsTNTfXXO3A7gIM7FTNyzvbptNJePRjN23d
CL+gByJanJA6SfsAMutmLfIV2RuOXy7oabcjHqsRGZv9je7AlJCXqbkPTREnMTsfduZb6epwgQEr
n7t+kY0aH/KSNQIa9A4nqA2GrBXP0olKScY8Wmrd7IjFnnGhYKA4RQ6wH0gUYfBNhHe/b/YLVEfo
tXbxhe+H7MfNAy062fMprPUKIccbMXoglb233132Z4B3qxwtIosYIHjrHK4PwdxTwSgE5BH+efim
WRKqVgwWliPNnu65jWcXnyo6o0sNomzUFVTvzsuJBL7QSjXx0g2uOS7FYBeahFfkvIS8rPTMFXog
bFPZfh3xo1AKrRtJDQfpVNhXpzGMH8g40Ixi2CtOd8BfKH1dKC2G/SW6n/BK0YsZk2ew92Ytknd6
0R4CPLhNzrj21t1JNKEuEzphp6ChBAfnLFXmLDXT5rGB6RRpMJn/9r22lhe8xSgm93rsBRMtPZPw
RGFIQGkD45JRjc4k+kktcS8Unto6nhCFbDnzr7SrCxSPp9w6IjEcbKLdbi4eybKEpCPBMG08Hp/E
nOydDZvsfJVdFZqC19RCIYU5F6fETxi/HFnGkcM5uKDp7lIUH6VcZAwSfRCeP/9kMdnJ8QnmcOZO
2VaY5ALmRP6CbH8+5NrnjmhYqxjCGQ0b0y6Cwpu5L2CY/EmNzaROaer8L6+sHsL/GIqYGugqLQCG
nbGnUU9E39pxc/Yc3NHV/uPqhSiDzXNNHW0N/rPGr9D0kwqveaqoUTAOpPNGK2GeXbTVgYI81apg
c2xuLLDsM0dWPoMMmlgIhPPuRkmzUhS/7Q1gvr9d2iP4Qtu+OLfmaL/vfcRNO7GHacp+EvWBXy9X
z6fcbDNM6761WNU/euSIqXvp5zg6vhYgqUS7hJU1dsW8ObuZ+B2jr9ggsGlwNFQcoXTfJqn7xgTp
h5SLPjc4D9u0RiEEQmr3DVaJElG+ZlpdPDSC4kyWXjVgE3328nX/2ukFYB1NJ+w1EZJoz2cLAC9z
tUKPAzOBwkoIA8ceDembL8jSL7PgPj7HZS+7WsA/o+SC6pRsd64jFtrsyz47W4hf3Xba4FElQv3r
FaKYsUcXZBRdhebPVWDH5j0daEGWGJauzotzpMgmgz2/cyS5aHEMs4L8lXiF+Mg896J8e1dXErVH
dvs0bDQY872xKlBj7ajr2XZndfiYsbKA+tlf+t4GkTsUv5djjlg57PMVd5tyFEY0nlBiWNHlbrSZ
gWZ8jmM9iKeHzO8fJZ0tzLMDLtxdWhrSHj18sN/BSuLuj0jT2h7DzVvkhft96+g1Z+LgVYxnE/WY
wPqyQ2UvG02F6diqiA5vb7RggB2MDvubrMOrwXs1sh/uMkQhs6GFMYk0oJsWC8chW/fvsu/Kp7Ni
oUVSV3CEpM7VXTVL5Pt6l2SCD6U5qWM7h1jVeU/QY9OHAjWDQnJPTN6aQcz6kNSsa0oTS164EyKP
YVdDF65/tcCfHlfaiFNgsEy+eA1MKXodHwGNgeLNeQ4Iqts6mUDGxcXEzG45AjejY0OyFpRdyBFp
H71sRV9YDFMVcIU88cf1gAD977xU6iOo65+/AcUsO2qOXqBSyKgdtl46fCTeHpTDO30EE+TgYdbG
O2VUtbda3+pWbSWuHz2v3EOtzekwCtd0H9rdYICkRhOSPzN06ugXUETcFpzpbbTLZRwK/mMj8Lo+
ddDku1sN6VzvR+MV+AN9VZqIS6zkV8da2N3v8VBq2VFY7rXvSfbs2FgXTu0YCmzxjVP0wvSuLRrJ
rgWEOZgp861Skyxlcxb4SMDBfqWgJiHtpmLyqzqc0Ayn7zRQfD1P17ShVrxWSvpkmj6HOtvnP+Mv
myAtr41cr6xC3W/RqiJyD/nwbrybKsXDxE6ecFv0X5R21tiYq44zk/o11jDeCiiUAZRf7p8tAus6
pbjdIqVDKG9xslzWyxoSweAhVSE/zpzb6mlq/KrONymrWlp7G6IhFFN5SsTXFj8fEx3b1WkvXpL4
vJi/w8D2lvfC7AXuEhG8jK5FQ8U9PkhUd5xvWjQcPtUc3N1Fqc6FKoElFBwpoYyHho0U2gFBbqSI
koHAv8C9KRvp/bcyt4lh1hYD2Yrd+TvTOOw9q+7Ggc3xfxLKzQ5uwfiuY6fKH2hgQqMlfh0kXqbi
/KHZoicgoWWkvfpLlWC3BUI4Lu63i/1MjuzvFwUmFivB9E6gHMkGyCUbO0H0dmRvUC8gC5Xdr0TP
2NRhiMUGVIYmVUcOZJLn3uLUfm5Uay0QEpCGcapU5jE2A2XL6tblVrEyoIK/Nq5ttUyPLPUv5/Gb
9g++ddEpvbi9dVdikgK9Vey9SyLdtt0m/uiqKbXK0UE9V+jQvWctN3bpTYs/7nNoS2O4FtoF1qPN
hwUzhTK9JmAgKVSDt6VzhdywwOeK1BhdwoCl61h053MtMNSWeyRjr3Zke/76GagHuFLF/7u/hT8r
40IFvMLBJHaKoUNe25GY7pzv8dRBZEVzEkvt3Gy2WQ1ddnId8KRalBHjwRsVWnZ678f0PZVgyGHV
szifX7fox9FfD8eiVBEPF06YXAytXAkilt2FAGpIbe0w7SHEt6KaFIoOIXbzYmzqppEL4GuJXJAt
tBBP4b+sqAGTc5CMgacBr78+oh9Y/2XUNPZEg4AxqUr4tCrWZDLYVVEyn75kT8kj+G9SSgxVG92w
dE30xQI7Scbds4G08RXwm+IPnZprIVBwjc2oL52TQh02CzhPvcRcZllWp9PcJYBlyhjRejRkEnGK
D/YuhviCfTNSZO2VPZTreT/aXnlk8GiHHqrn1ldwzrtzoewnsBALVvivOdLkeKxl8aW5IxuhLTeD
oroiQ8Oqt3KQs9dspgg0dES2OWUbSsb+aeGyIXz0n/QzPvgSd9rNs9zMwTjzbadTzGjncehWpTOS
Wm+0OSHuVYHoWqLeIKC9b5n83gIb2ZEWbbTMjqBmjfr4NPV0CuxpXyCPt3Qtu8G6UMHkRhuNgw9l
WDlePeefxnZbQw/jUcBfZgCDlFed329q1J4Bkqpof25Ydaf+5AlCgMVYQBWwlFNOib3ea1OpOc4N
NxhMj7EkwJQB5cPoj8ySdQ2ugDOUhfUfCNCXZIKaRBVfymyr88PDDgp9R1SrR8D6RYRBw1FNY4xK
zX5UOdVcg8WEg+XHv+Svx2wDZ3POpltMWXcKTwl/f/JY3UFAY1b+BHpUlnXdlMM7SZXdT77f2D0B
4QIuiCbcayefDf48uHg5znsqAxfLDFlM1nFDv6uK8n4R/tPFOaeukEzuRxHAPnJkV0xGV8acaX6o
woTfIhcCunpHP5HzsYOFtv0vh4iDKlwn1DIQP3L6EJaRiX4klKxnYnbQUXp6hKqC8JhcFY5hx18x
FaYBOUaPfRmLE+14+gkNV7FCseI9sUjzXH+Vm6+IFXEqRt8hvJ7uxrcC9wf3vSjeBB1sR6k69S+j
ztQMGjJ3yd8M+ll7QVeGeXaf0lnQNaxD4mRKGu8DJWkiTnkdcSOOmiqi+QjWVd22n0KrgwL0TM0G
Usp5GUPelUkIoll4qlXPohY8kzvoAORXq1nwNFXcKYU+wlEjwxjoH9B/xegTB9Qrg1OMXMDwzp+q
IJJ5NE93tAnKnt9WVZBDexh+ewuHU9Q2vR3nXbYdzUyh54dFgXgB3vzJeEkb/9BywKTmKxMOg7oQ
G78Ms6M6tOU9HAJUOqZ1OWmofFnoEs9E18hMr8Di8+gud7/y+oJ/AluC00G1qhZ11yGcDLlPJsU0
sK0JDr4Ur6j5ApWktulnhxLpeaQNJwsiIzTzO72aA9pUEkiPpUnfCoi7ig1Dol1srkvEuuIhbprM
/AhIpe7y4HeMo7xmyt5IWUiGmC/w4GCAjmOgPGnveDp4agFvVN94BAUD3+FmyG7PecqUZmxPs3DP
T6kgv6U3hqgWfMqe6msYl9ViHfnHeiJYEKfmK86ZuiK2xAagAnCRB7AKUa7buvZjtiJSwKn0lDbA
D79mdVHo06qYyXPPF6nFh195bz9oG5EIzcBjcH29S0qfCbiza5Jf2COEZ4BwRUUn9iqQZ2dQPrBM
nWfU7CftUCQumXqkIiPPnW47KgPDlt8FSzbcbOSYPBX2wTbrlhkw9kcWhui23+pN+tB3GMi9sq6K
+x5C1hCHSM/aNpj573BdKs+moT/EwrlMv9nelSepCQxRYF8VV3Rk8jHSsU29ImSjFyOYxxgIiT8j
IFLq/f5cXUZYKKH53WUkC+523bCMFH9q4NQICBpuQRV2GczMK3TvDqY8VH/35iNPhx4FyPFOKBGc
SlmGd93FF6fvr2u5EC+08JZQlSL0uwsvolkOriMuu/S+16m4w1M+rLoGk2hGijUEH22J5CgQLfsi
OYAm/Xpo9nb6vu2GyCA9TtBpL1+W3I+OqRqD2ssfa/o4+7qcdORicBzZnZ2DuldDR8Vmi5bDQI1G
ERlb2hebFCitmVYtdv1wuQggUcLQc1uWuT7Fy7TW0MsVh5Gh23/IexZVyEUzqYz6KXTRZYN+v/1o
M6SLlM+EzZEsurCfkteElqlVDKbTrRd1mR5yW9cbW7xE/vhpnn2SgytV7m1zvPClHh2NaQkIqk9f
HEDEs9XonP3fH6rVUzkEtLU4e3Qe8hXQEO7Gk4tqFBStL2wzzvE/hYadl2cSl7+ipGQJzt+QHGqo
Sm72Xks2FOdH9i2JFe/A13bm4T8IDIf/LQpQy6YoJK06S3OlHTv17JCOs3rwRI2lhEtg5V3uCLEo
ZPQRAEqLQKqShmTQjoKChWtMjRuwAy6W4RJSJb3O1GoeVHmcJmUcftOBzS/WJnlP/KJZWjpH1p6x
9O/CRrc8w9WCf+wM/l2GnfmmWlaxufTeiXieQviYx4Abwpo0SFm/XYIk8TIbfne6tnlCh248Iyv7
uaYktMUhv0XKAw4fokXFqkomzGUheLN0NWwczbhHi8bkw0FCCY/K7ASSdYZrf7PuV9QueGOPzxzO
9Rvh8QNGDjJsAcrfUtzxcnLIfQgCriSrqKJfQO2ZGw/KSW8KtTgvtORPp6bFxtfG4cnSbUeWDTTL
5G+K8996X7U0K0um0Wu3pDH9qa3sfOp/inpPr9thN9d2yEvKaAd1nuO1G5CzlsbVVovxBRKRGtye
RFnEOW0uZ3DeqSX+CWLA6RhPBqNpfF/6nVomRzh1n2UkFvOUq87BvtiG95mKYqRvsFORxvHBks0N
Ll0gPNyTyKX2vtIMruRFmyXxMWmrxjkK/z/Tyc7FKUoWE1KfR3P1HxqtkalWVW56w3OrkawKhSGY
f/6fP8uZU2YyWPubL8bYtEIlO00TG7P2dR+PLTt9xpGE1zNhQMWY2g//xLL8wTJ+HhTwVBhpF5Bn
aEFNo0yPaC9SZ1QNpc25jeAlziZDdqHuMoQWXMjsdepXqM5cm0nYMZcoZqqFg9iJXkFCQwUqOgy4
IrzBQm4NGX007v/I9QqBAC8D9434uq99SoeLGEacK+j8AsdWAhWj5b2VVna6imoAMxnBrqaVRgkX
60IJGP5wiszOrHnCzk6RDGsiM6fACBJ+5IMCnXToh4k+AEIg6utr6nlGLOjipIB4TLuvPBXSaT71
ZAIoGoNRsjYSUmoxRe3YjE9P6DreyAOVebqZ53xqodCE70AmrVC2I+Ry97OOHD3wjm0qBxW9x0In
CIE78yKfrjW2sondX2P6O3oW+rW9OmjZKKw2ndpeBelah/ptJtd374FEiXBuwfD9mzRAON3h59YO
iEi2TxFFSuOLZb6ceS8YrJ3OeXxSGkChw6DbeblJLj5EbTjvHu2gwuYo1FrhZB+sadejxLz5cUoZ
XQy1vpMnJ9sEPorakcjtcevUExaCp18GP6ICErAdS7ueu2/KCFrdVSyoLzQWqo2gMKFL5YEpDRKN
YVBuR0sZAO1V0fRV+D3slboXBI5m6KgLSe/2d/D+F0PF7DL5JANhuR/u3sMiCb4HOUYrXah5/GUl
EICtRw1NItAc+6mjWKEUlUjiRVANNBSNq3bk6vd5dr1NPEgpO75d4kMIJNFvt/OR1yRH1MlwzX6M
ZbS8zO7uYL57ni4UchQe47LIBcq4FrGYr2UnyrB1JuQmQnAYGKKono8CUftaYxTwO9Wq46fB/2nB
UqsehaLRHt2bX3O4nKbOWRHi9ZG7yfneXT2QvEmgGYJYDR5ae9r7BIStubqt+n1C67ZUjRg3OLKU
BKffq9nZKllNiFBw1BSXhK6qdr5Tep6luElKc/6oC5jewLafgYR2VpIqO8zvAelSTNDHMVJGW0mP
MQJN0SVUE/sVFMAyVnyOWCgVwGWelvXVw1DkX4EnLn4ALyWZHi9yt18MuJTZXbU9hW5H5U/0wAB+
Z05Lo+D9XOZXAzBhWarVaXeIQ8h8FrnEhiPY+3/SiM5wkzpvnLW7nqCkwo/zaYLLNGEhc89I/zDi
/siuFJDlBvjt1985d/pUNKM5kVdkW0uC4cAyN7HTIWLYN3bMU6SQkK8/I1eSFMzQ2DfMCzcDIdoP
jt6Jg4KL50WwM4unP2aqvHxokUyKHobAd6rp25lOZYFYa4TrAlOrjqGWvRfcbOe02heitSPw5aKP
p131WBjmC99XxvbaYqIHC5Lmy4gUGh5VAJvSizscI0qxU6zg4H+bjf/4cV6H8CI6OQPXM8kXplKi
Q3Y+Kz0pDXu9zYCM0g+F+ChZTK/kyX22YVfy7Tu/Qy/RN7kPmGkmnl0/Ce4jeXBY/nhwWX3SC/mc
deCFn/wZg/F665slgq2PRkMfsqLf0MSWuS2yCYeD0duVHSkyW81/1EhVGxhP9eXDMpq63SkxlZjB
8WVspOQyr17FxKSfbJGy5aLl+gSd5v8Z5dID2wzWevhtJCbBJqZMxCivKR+EhC8rhu+pgyH6eiEW
zRlw8t7sJTbjmNIBMcZbYTVQBXXcZw1iArhX61Lx4mVbsjdCYQJFelC5B++UzfLhK6C73LT+Xlm+
27HdSRrywRNJyPz7g9Z/duedE5P83JgaOzcuoVlwi1B7D8JmnWdtbOm1aj7SSC+DVJdo7mFdhlgf
MqPdXoziw/2WmTPbUVeeyTdgDMCIsC2XcAzHNQoxQvNNYGEMmWxTWFBylFP1AmQtLTP/5vin8eZB
xUUV3qSqN9jEonw2DXpIdMsXfdMKMw509EmqFDco1m/Vtx0Op9Cjun2bVWJnuJaDL0sUCNNHhr+x
ma6FwKAObc1Kw9Y6pFjA7fkHa1FmGIYTIvxf3EW0tr2qSljORURyuldx2rFUMqGjKOWrYVksMcE5
jyE1PEdEz42+ZkNDGWZPB2yQvHdQafRJMn1t/JbkAoAt5UhO6cetlLdQGSk9cYHI2LI/3K4xHEg7
JQQnYFI12GyMl5/m/pu8AOd/XB0SKJYrzsAaXVOTS1HkqBMB9RBRgl5SObEiksdttVU2gOOYmoas
vhj8reiAr6SZmh+3gDxm1qm+4mO2A+layIKMNY/XRmAcFY1Fltp31PyF86rH86cItFAHNe20+VzC
IsvPtPN5Sh3wRrOKSQ8xZqyXeySjVPqwqJigwlWkWkTa2d74yrRVed/lr37ksQAipWcCYS0AO/h5
QirZfP9yFFY7mS9qcLmhQuLIoOdlIG2uh+KGz5PFSaDcnYwAinQI0GfTD4P3R/V+eQdGkoGNoEZo
eZM1U69xbZf0tZVS99+HynZaqgMttKa9+Imw0x0r5Pf8neh+L/PsffvUPmFIAOHNpY7O6JR+bC5N
u+vnu/J+cTVQumauP0W5yaiGsGHv/gGgoxEN89jKPQfOHNzMKdG8AbFRH8MgG9YlKcX1PkGKdHNd
gjRixQCE5MC5su0wOFQVZoaD5nebtsb3XXb2PGj20LZBC6VdYJCKJdxNJzdudqBmfhmSEDKWdoJw
zPQK2ZZPfd0moos9kYHHZesKfWhC6N8TO4LmKTl6kDhV/5lAVTM2PhsPg9RhaqqcYs4kHhUNTnvT
FXjBdgX3Wdr/zaOG7NS1JFgqJmQYC5S27hGogLBWey9DnsUjd+9zVFV8NNpqLynI6xS3Wqbn5XW0
5RFfCHMeV/o/IenPxYrMdhfdbSy637L3fDNGwuxpNoDm/ZfAX8FXSIjg9y5UrZ9aUP5QtRo4H75I
pzp4+wLW9B0TeuUi9OHVg9Myf4V7TNVaHS8cO+bO7ZOno7qaLH/HTps9wQuGrWc+uv8cgqwGwk8Y
mvjTkPlBigQNiIVcufRh+m09nVIRZI21ObpTjoqafE9aagLNR7fuhvmC1Zwg+ED3ynyaTdJc4Vjm
OD0HTMxJARtzqeDgmkEGyctFEus5F4ENJlbwA8Xz9UiS3EdDj0PT9BTufBA2ENihXuWCWIWamuJt
kQ5qfxUcyWCxh6O8yqM/a7ci9FnxG4vuoOC0lyCOM+C81v0oJ5on8gxkUEMkZKFe59mZur/Xfsx8
JGdm1ODNIYXfvrqtCJN1ARvpW2vBhfmBovay+ik7eDbVpHm53Me4FPb2uNf2vKcK9Yi9ES4f+6nB
PqHdhj/nTupS1qukw/MFREOophKgTb2tpDZQqzvWS764CnXc3Cv85BwVlpq9KaToZ3YWL4i2gWvF
LvsIPaRbqmX3cZccbgBL99q8EMu0UhaD8d0pkZAre5utCXXZGEt9//J5UpLjol+dECk4GeyDFFQM
S79+9C41MV1xAVZwklqy0Aj8m+15Z5vrCeceVgSUmdS5vXj1MI2ZW0x7Lz4FqZ/VbwUFMQlE9AMM
yeLFdkxiUN4pRmjyuKngeLekt3gLBr5+CaaFc0SkuOv/01LbUFD1QOkjCqs1AQc+S9rwotvFH9UZ
NHHm3X4u6m5CcsKzrxTfxJvz7fTckoBkIUXafUjqNFMg9wjwoHJCT3S6T0VPrYMgQMd/edkPTRE1
9K3oonQtTzguAIG2W2v5ssU5wwhwaUkBz5SIsSn6NObwnX+NMlG5ygYL+MnKmyNmEUupEQyb0FCJ
RvimSMIIMO3UHz2upsQa+rj7BAStKN3M01nkzcz9IovA1Wur3/rm2Vya5e+x1V6s+RfAaT4fC1RP
faqnR+dzgTsegUs11+BLc+yLXbzhOdjyBdQVtX6oT/jcbR4j+ZP2TXywqS0sUq0YIabiEo98O7Lw
ILX2clb7UZGPtzA+svVlU2a+QxXcZ1PDcxotBEkyclBwHLPtuA5XcBXpgt24f03nr2WLSQqmX1P6
el7y65wBMHPrUoCoeNt24yzP1W5zA8Jo5eb3TYha4UEYQgMBlrxj4G9ke+yQ6kg4RqITj7zNaPwf
+ynZRSQKdGLn9d1/Jt6ZokaWmD7gmN0EkQ1m5RQv7KO2oo9zRjQKldSjmW8PtFEagswdlzfiWyS5
1wJjJhk5yoB8oD2ob3j19h4AudojTcFT8YhizYm5qobHbOzblVVHVsx/9bbWrSZR5IixTLkIzsXD
5bsW97384bM9jLgW9JbYfo992hjB2V2qWfHOZV7e3Nf0wxsyeWxbMLYldAcH6MOvaOWUvVeyueK6
xNyQ8NUcajnV0l1oUhgKXBFYH+9dNj4HbYGuPytALy/JMfRFXduDO8Ab+RtFe7/mZdtF6zDp5OjK
2XKOW4IhQTGpIw2NB55HaGVth49PTfUUk//chRKVcnj5pBW1Nz8uESPeG4Jz5hVIT6S9/YoT9phE
Ov1ye7DlPkkpsx3xY+KbYQiDZHy2Ghf+3eKaGULWp7Kh5u9xE33QOSVg1BuYh3XMHEuI0S/JQ9ZY
wNYzMvsWPTZCMyCNpwGD9mdmqXV8gICWloFKkR8lHmhqrabMjXfjp4TN03jWn2Jsgi/gXZhJHJle
vq56rGlTzrIS03ZdAkWg01OqdJrrdVr9zWDyoluT4n9joXESyQEe55okPJhXsCMT4T3E/MMglM3S
1ZByDM4bf51A5g0WyKLNiOSCT3sCKTBaJvOKwJVmYCZQI/Jeq9q2qyiAnX+69T4q3OLobTVn/jT8
mn8hpPSaknigbLnPnDGblESUDN1hSqPyaVHPwISTpruCAb5IqGVoG0HHWLgvGKQ+YLf3kb7lH/mS
bw0fK52WuEIlRcRN4CxMMtzo9RRpTZ/Hxxn7W63+R8IfaddQI6RdhWt4/IE34BL5ZO0iIEhzNSpQ
RlLOw0iy6P4yLa2/e0YJeytwxI0JIIttPdciBqM04vudnmflb3NFaU2pgVW3XSmNKGnx/GYL/avp
tdA9PiTdksl4yjXRigqn0KepadTP5N9aFAB1irVaLbD84vjsejnESsHs0rHcxZJYnPHbpBFR19OS
XmXfmkP5gS5DaO9CTVETUvLMHkkVcR6/S8aGQjadj7aGG+BikMTbdE+BenOs2SL8S2KDeuFS1EJP
Y0In873jDEhURRJOJrpZfWuQGz9jaiMdYLpieHevLraItOKI2rR5iVDZ8e9OVFLh7quGQ6p5YBQE
JpItwDN3Ok0WI/0ZaEl3bxLM/lqxUSsa+OmsDe/XU7q2qxkcg2D5LfBTd898ZMRHJnjSu2Vcyc0T
SNN55dPJ37sWGpvblTYnwT8nGdLtKkHgI8CE6Y7az1Q+FUAJPMLqXuVhROLWbxvIqtgEouqjdFsK
o9dS72KrR1W9L6ktEPFE9hUmyZdtda/66kKCnl0m9z6Nsi+pZDqLRWahO8j0p+RjDeU6kjXZYZdv
CApRsg8S0G/RdhqLHFkDoSVgAoITXybXJxcEJfi2U0oWw4AtAcWy4QPcPCL6LBFF0p9eQxvzAxdl
YV8oN90V2Wp9vjEl6/W0zxRUy/A05DpIjqOmhWfzsp9fXQXhoQPBusjDRN5GC3uCXdKBO3QFAUI0
v/jEGdfofvq3wmxHkq37c4UERDRrFPESmY+yMZkaqlo0wU0KL3riXQNF9EtUDhp+rdZBGHF0cZOj
lcxw8T7kC/gpPuK0yiRvqzTd5JiOWj0tmqUSzmwmzfnEY08UDOMzbGOY+se+5iFYv3GvLiXAREDu
6l1QFVw0RSBY/uzm8ASDKb5aPiQp1JUq9cervsrALMMw4U/zAUkixkoW7skQbiXZy/52lKu3qS4x
c+Uj2iAvDwAh7dU4Ng36DWT74JZ3y90HAYn8Vh1XbWGMrdcyJy+HCkDKWKc87bL6y2n002oxBb66
zpmII/5Jk5VnTMUOCs5yprg0SkVhcEUlowubStDW6J+aR4rKdp7wwFoZdqpLIT9IM/utiINyZmrg
R63Ug5PIlyVLIsPkzIj4f5g9oCheQpM3PwI/iTZNPFki/XCPQ7WmWep8kGqKI9ja2VAs4+aCh1UJ
SSi+RDOvPdabYubVoUVLugoXfU5Av8bFx15jHESuSVD0ouL5Hufv/7cFj6+5oo5dHJLZIYfZssUe
y6+D1Puva05s+x5fpCJTd1MS/kFopssrcKDs/v5kwI4ZeNE4TVPB1usFOpScoK5HmDgG8k5CiUfV
Eqic+elf2F66VyEpMM2YgsAcmNEgIr3dWWsFKuxWAw/FWGhcJOOU0dF1FznujrQ5Evvg3drQ4/Mm
OkDIyW7LXKIBYOxeIdiOPQI5LZ9XsyJxpi5V9k6ihMvsFNYX8RZslNcbfcQ5EkfcXGSfyvECTFSj
KhNlBfgxVM5epETDHA2D3QyQTelSSyFD3fCzYCKJZ8n2Z9MmyMpicRdPv/mNNzHO3ZJ7GFjsIJPy
C9QeA2ze8fZTyaF+7gHjhYuVbHqSMvLNWkhAh+hQYiDYiJXUXlT0rk+bZhTVrt6dsYzhNQ+f2Bzx
8OWrorXVlG9Uv5x8UShNR8WgTEaC1vk6CXNqCUk/7s14y0eoutxd6Omck6+i4INMwYb685/fIXT+
UnCpkgLuLx5I0dkd8044VDYc/rapBbrT7l7XD1lBTVZ2Oq/0ERJJQfTRqisX+WkPjjwzsyVvhaOF
oqThkngMSD/KMCGaOSnKTWPynd0eXJpZithpsDXNGiQsb9c5tkUa4FKlje3KB3x5IcutHKpXpgAb
GawlqzAW5wlv/vtQtDVx0CAgrmwyvr9OLsHaT2A/B+nJoqD+NTfq57a7AvNO+g3wwwp9yb+HEWME
mrG86NLP90tLohXWCfFSqUZNnCPCYE0qVeejhzQrSPfb3AbE3K1OJGjy9c3wHuAZlTgE2fA16ejl
T1cx9W+xqKtIIiJ0Q1rb3tt9gKqhU/GTDr3SmyBo/kpZYb5Pej3QJeP30S++Bvh30dU1+wrbVBYU
uPFSXQk/0af0N5uAHGiwFocsxz7Yi/4wyMxz5F9nH/fMXDS9kbqLHUyslZrS0z08JGW2/NsQloPL
kymlPmbJ9Fp2eMOp/fXoG6IP100yYNuFqT3NqOc3xj3zlq2Go8yZUBnPK+1+wvGyLwx3MCujC8X9
snRRY6HvBta2zLOHCTGRpOuYEaxZyw22wvUdWDVWubM9duKeCmABiFnLxJQ9MBq8lp7QUllK1XXo
Y0uGp3BJxLRhEgxK9ZAvqhKjniwAELzKJlyrOUMCvSAOYrAndkPBLzpJJ+6IrOGs5YPMQLX0Uog1
Y5GSu/KhDa/A6FaIkwxgtUJ9rOQchUeEWEWRz1Uam5i+pAQ+3lGjLKeHqvrJ9YBhLNLsiMYZ1UOl
5dJOEUsKpEbmYx0wq8CfS53EXyyfSj+NF5kteag55OzMymVx8RDgnDZyLZlA5j6u9T2Y+Rg/2+Vn
xElgM0zpVNubFk6a/+7rPsQUoewUdKCx/yCVvDeSaWcb8rfm8iBnAH2y62abTuR7n9BTy+YFmGYA
LoZoNPKSPhbW2G7uvYjUmxmKm2nCmz+9JIbiA7xGGzFCALif+fz0lA1+4e94OCK3Uu2XTcWptJGW
MOeEtwtVf4xL4Z6DgLCokWAC0WA5oCCR3XrVJerinG+T0Dyt97NfTRf3Yw3h5vqShCCa/iLv/Y69
xqso1iuuDsNmiGEWN1oNTWIDJNRU4GxYPxozv4nTlbr93uDWXZEkeBf0MPLHDkKPHM0ZELIsD/J+
0z7QiFley8YQIkoUXJusVtxOFL2sWmLmdhp8hApEtgzXghJOgFQc0pVS8MVcmrQy7SdoNa1GNg6b
zRoOJ6+WTwRJutTsEPQRa/dVRNRMvNEC+5yy2EC7JfgIwas3p6hELZ4z+sFjRQNqDfiyseF+CTtY
PU1ZQlKF6XCKFLiYPn518mvEud9HvG7cRTK6+oZOOkTo0gSr0855NUoXionnOgxdZgoJUfOmh9Lh
ic+mXir59+6eXV0nssinK/OJpbFrs6T6IDFNTzJgLzccXlf+u9FrYsNA4buMRWsR8ncsnIJl+wMQ
0EWbPGoMMLP3y0PyTYgKRiOWgTChJCRXmCSuCSbrthWg+0rAEAlo0R5LkhnlCImzcve5noiAMFZC
wb277IBC4fNeuzhtAH/0b1d9+szLnwy3I282bUWWh8OUAVaXjJRFHC6tDcwRbH+3iDi+yTsbrZ2Z
lSH9UHv1w/Ok1odcOOeBNgaMj0m8TfzUNUPZZ0AWuRzEcaAlgzAeFZmrqsKC3bqr4yWhc4cQV7B+
hYoa6UfTBlYSNSn4KGYBN2aag6G5wEKv9ognQlXk1Y3MCQQk5TEYBBBrZaxBtkyimScS5xZQSASi
vnyYedadS7rkwcLHhR/mOtACGWg1ZnNscKgA+ybrUXlALriYNcedtyuUVBkZNpFyIZ/qtk3xqqER
OzzoYOwJhnkSu4RXdXDBZcnmbkMb8QT6mzNdeWCbIGSgoDQD7bvMVr49Z2JDwdpMUfLbjIgvRIqO
CgxwLW8iUEdO53iiGEEVNtnd86YL43P3w/YKqrhK9X69aTVjNKnG8W0oWAam9ST5YJrzjbZUYfIG
yRaOcF5JtSO6U4rPQD5+hgEegljwqv3hMiMY2acp3yqAxPiCgHT5qagT4Kn/JVoptEdP5jQB3Z2R
a25zKoP+yU0bbis9ln/J5TdJrUGP8OgfU7b913bOYG1PJiYLs7YmJYxJdhg7muTRvkTF1BS5E6ld
IhgMwhMB1w+3myw76Na/CqHmndu71GW/R/8osBthNp0YTjxxLXrAq+l3Z5jag0w6yCogE/0prV4v
1feElXWS8W5tYoYQiHgmYwcpJe7GFF2fzdbnPu27QAJzzPb2R47ZomVOKV06/ESDnm1AB0n//CxM
jtj7wZHy98TmUgA0VRxer1mD/S85b+aSqGjgeEe+4QyQ1Ahpqjas9bjbci/mTRR0KmsZLDiuYgdN
U1V+r/tASFHxwX2AHr8iNVuuAEDUGZc9cjUfHjHxvw/gfrBG6a4jgtgVNQAXcQ+VjDxwAwIpqlCT
k317MUR+IxA3jhzg0XMrpLNDBE10WheTYy4M2Dpj0sKFmxO73cgSKDni6cQxMwys9yVYGK58QpnF
UlEEqzMKxXfqqGFHINcPKcezazaayTriCoJmOpzHq/CyzaLuJCu30nLfLyQ0yK0q6lzlrHAfqroT
9K82Ae9RYqxMODHPkDiRslY/swMxNKEZuWYFcjzKm0Cx5J22P3dDUwz8gpa9WcE27NLA08Dfe9yt
CrteEx8X4/eTjdCDGNzhfqfMexOCYsp2bVQ2AQN9F6jL8oxKe80RCAjyBmy65qCZLdNzbCZ6wwPc
D/LJAb0xPnz0R/0Ev05XlelM0nMJIxGLyv67FMer1tl9wn1ypYgx31D6tj6G8kJlzzyXHIw4llBz
SbjNLjj24dfqJnqQ+cP6HF6dB/HH0TE5JUJZ1PKzPwsYm5XnbmsTXvBs1J7d0SBAT2sy5LO3CyPo
iXKO82VUtaEIwg5+t4+dWsEi1arlBqkaRcQbSMs4YD/8AcOwjwB/I1UjitJh3T2/9XLgeO2HKKwR
ZIbOYvKgU60hJed7V2bYTTNkNHz4ff0sKjfI7h8JnoOXl2YrdOE3ndd9n9F/r03NPSqiUdr4W8Qy
DZdJXiNJlpjZihfYIlPcEDm+Ceonvn3TE/0JW5C0J14kFXjqXsqwHcQfdz5EMZBF1vZzb6yn2d0C
pA5KHwAgZiL4nZQg8lfEGL2mPLtadEmyZxv77kD9kX2+H5ooTt9IeKrRYXDM+0dLotxCVPwac4Tv
/0bJzZIWhIo5o+6FcYMf2kwbVAIh7Bn/1C7PE7YPCAiZnaxf2vINHdFIf5VAP1misxYY8Es7/HU2
TYDMF0hx07vJ0WdDuqj3GYjou+vU1nih+KEh9MgtyTWpuCBeVWzdnBMWsza0ljO/Sgz/PshsTGOs
ZaABTKhbvFN2PhoWoAYTdrdlh6hxO6hw8HUD4wtKNr62ImOIzCP+sGbF9iH0G0YhccuGCG/LYIKY
ABvm5TmauYPO3/7f2IqcRok2QfsH3kdZqMcyESIScjfoeDQmav2AU4RVxpQP2ZQIFZliI6YXs75X
T43YRdSbzL1/BAA3doVzsrOItPXcjIRjByKfEOxfRd0DhhpeC5EinZIAoHqfrXCxOpsbAUbxNWql
4ndZgRv5atm1a9joa/CQRstmt0pWvhf+0Liq0BSdQObZQ9iq9+Q3vSnd33kVHcrumALJ0PAGR49v
yyl8tcX6ebMyRPWPp4xsoQK5wg0XaF1wveekzEF3xi6CS+dtCh1lkK0he+eOFs+VJMQKmvXE4e0O
bkhpJiPRKi7KQ3UvGEOXlsCzVxOc3LkVp2bc8T8GDVxLmR67ZilwWgh/MwEgj9Q3EewX1SADM1HI
UqmX9HRH77U4Ujo4aXUxrnU/FLs5Y0DphZBB0uvrtunwG12lYkYKZQVA++tRtl//JL+w6HmxOBHI
31zwE4ss2XJoSM3NoBThRGd/zqvBUfh/K9kN2gw6jsZeIFuJyRQYGKEVHvMqZ83ISsiOl3SjMKZq
cuzbip/5QZTNontUSypalWvMqDafijnhFsrOGRQFDXemtlqv4JnRo5khbTf+uIQ4bo2Qq2y8HSGK
ocWFcCnyVx4FmSsMGXFZKE9vlaMYf4EYzkOq1b9vvq4yKg1GEoclDhWtVHIGukvaW0P/IAo3WScy
9jgkFpDGppU7f0hBzpzLBbRKR9IiVA9R1XunoDICMkxfC+QABw/JHXXEMp58NMK8EjTazB7wSJrO
q5kiWoyrdVCMf0nNVFfftxqu91/ihibTX3/9A6dwfCY+kAfNU67ruXmpXkqjKGz1CWCPQG+uwcRP
nH3qRNne0nLofpgckmoOnXJCIWCtBoKueom3RF/vdK62r4buukBerGaaY1HI/8qhkz8GdmUjX7XY
2cM4TpXCZcesHrp27EGmnG2+s0O1iRha40VlqrSmgtjyrIDp/DZ7ZaSiPz6MLDvIgh9OyQEauilN
agu2q4zb7ThOO7LPy1IKnQQfHXW9SuXUU4J/9rRMLvuq0DgHK3ugBnnOaqsL9iBSx14IpJia1Oha
G+9HjAncLClMuFs2lDnOYzjR+5xfzYwMD50sx40y3o4x71O4RNC3kh9tn7J8kDHsQ5jVNpTgr5eR
6hmRdAROnz0GP/zj+kIUtIM32rbBXsuxSkn8WffxULU1GjlR7s02vevsCPrlLxuiy+5UxYuRe5y0
kHxHSoUFJYyCDYzl//uLOfzkta++MNu9JyMER8kU+9S/MbU5pUEN01mvzM98al7roVI9SpbADieB
l58zMsWuBEN4Ew6KIO1cYF26tsfKQGaWO9qa4oiSqeO6ob/Hsbks0bbTAxZJ+6IRgvaEEa0aFXo3
V99+fiUD0Nf0O3FoajASAAunuSfoybs13zhzlGg7w/it2R5CcL6hGvegk8LeGsygSBynEWhiwWOu
0w5ULoaYQfGk9ahIJARzCKLRh+fjrGWKSVa75CjwsKNQ+kz2P63Wg1KV92T6jVkDsnM2Bj6V/BvQ
VNs4m1QRROIcke0TAGPWp3yU4AGDI8uh9QE9Cj2h6vmHQiNqN7nYOHgFcKUkWv6apVIU/AmxevNm
M6hxWtPbL0w9VKDR9+0Z47cwq/CcR+9NoNoXNkma9uYArC8Iq4sm77j3MzDMiqgaE3tznZ15+OuW
51jR/syVHwgdfxAk4AjqZTZQngw4Hq/dcnMZdvXUT+iObL86R2ycC4IlrmPyPcW4kthReBnAIczY
/RAy1FjPMU9ZZe+MLS/LgNQoh0pmOn1fU9shLSuCoTkL7x6ThcZQYokyadf6zuCZVTjLb/AZEGgo
uEmH119csUu3lSTD0H27iEIbPePuUBqg5LAB4cRCUWEQaaw9KmJQTfBTNasQjcVAhepuvRxKwEB0
1BxGZZZtx/kq1zhtfA+ksp+fOyMiwiEpoiXwp3bgQW08lKFbJ9EKU2BA8CArTDsbyB3YMST3N82Q
zAVy7Y3vJ/J5W8ughHOuIJOc2t7Yl5Pp796z2SJHYiriNb0UPj/HB1ovQMM51d8E7H0oXqGnLrdX
NIcXA/ZoNDG2Q5KXkslRqdvToutw6rvxpWBURWWiaekMs4xazSOWTae5OhxtQhnxBSh96nGxKXq2
+geVTlDUQmdG4ecMTIFsuYyDN/4RJ0VPGHciicBBlxIKHFmtszk3FYBX650tb5gDP3/CqOkQQGYA
/K3L5pyPOlhYS12squyng7O+SBgpfcx7G99q2OMmRrg5rFC38QSvptHdY6zhydEJkGvbx0YJw854
btB+vLdPjmfkrOMd5EdQuw+kdvE0/+qW8FUZ/D54Tc69rhLli09mz/CjXJ1u4kDK2ZtI/abzY1hn
X3f711s6ngxb+Ci6HO92w0JeHX3K6R9evStCnvLcu+dREFYp67TRAUI6mdn20Y0ahSTvD9H2HHk2
YQTv+sz8BBZz9Qp1T3tLDoqj4VJXTTquEby08MUNVIEdTZz9Ku3YeWbCREESL5Z49rAaMcg3un5e
JmufaonRIScG9CCN1Jt83iJ74cdsnUJTqjlQ9RSfoBMlLNwvjmBvQfT2bvz5b0vrPDsjermx5KCL
HbXGZLJ0l6nX/g2K5+mp8N7A7b33zRTXd4Wfy2BiOH3zdxbDRCpqJGyBFegWgJqDiu4PaK8MSNlB
y9I+z4gwPaWuMNp7/cc+4WeHWPppczjhfEsa9Msu8rc/gwnGky919Ag+V3rMpkeGizBC+cXAuYDr
x7d+SMx63ZF7Vu+ZNZSx4SSEE+XerbDIkEW05qMVYkiNj/X/kDyZiLbrOo4K1iyLD9L7J4x0dCwS
3Ok6R949KvFkOpYFCKv1cLn08Yl+Px7WAMkUfHbl4nAWFihbTOUNDdIlz84Gx+NnD8bKnR4HSov8
uM5VfIqj2or9QEnZQbD33YF2y8vl7qqLz6YBqg3BO6Ysb4Ncpy+vGbBKfTM4sQqBYz/hr7Rz95eV
cu7Ykc0yRpqPyBBhH/7D6jhrHlcNvqVuL5M0gzJBi0FT0QHZMLVdr1Qsx9vGL2hNXqhXmNgE+1X0
ih3AjFL6O/C3qStIBTuWhmJ/XeTehpY9pyAWu1SV1bvAxjf7WnjJdzP378KdOiWoF07KPWy6FU8H
W0Ku3mxsxOSPNfzMSYrx+XL1aT2jIjBZoz088lIQs51NtjmsS4/vAlgEm7DR62Wl9jAUhdIBKe7S
MYJIyv1z6u3xm78N3U9wLmcv/eafZyDWEb3XCTe0Uds/NZ1LhTQIlquA6nAhPA5xswx1Fc44o1YR
cQkjqbB8WeQCVBgHrJJCPVg9tYk/yKul4sE+4iyWwsOgkW0nlJwgl9D5Xo6D+6IywVQLMlofWUxV
e63KavL/nyu02Iuv7aTqZbP1C3V0uzB1lwpamzK0LpgpCBlDlKjEbN9FR9k0iZFdlLzl6J+jaG09
HGiEzM4U1/j4A+tt6fnUK47Odh2vsCRdk/A+rtZZtthGtvo7hRRWArjhN62PjNIUKdrkadquEL7d
1xUMY15FnRzLA1lf6IZNboqvYjlGMsav01JasNR302xdnFMALPqJZsl4NKPwSiELQ4KTptGYG9n5
7PWO6dmnGg8JhBUoy3PvgfqTibz2MG54QGHd/L6DwG9CibKStoZwdE3Yov6WjO0x93KZPAJxjyd7
P/LqhABp2JEW1unnSNrfICennE7H+MmV4OnaZQOT0XNlCoZY2qGzMbzzsHxFlzIvFek/FCK0nrFm
vgbaKvgnMCe3L7VCLdVvSDiJOMBzyjlBsIzmz55enOvICwNuc9HZYYi3DApG7dQABvfMV2nAPbqr
ChzGcGgkeW6/3TxTbqsfkwFc6FVSFAzIo3J1GZjboyuPxbmffbyovvQNjsf8okm1ZXce1XQGydiQ
i2WfbjLWlc9l2oTCEAdTJakBYuJM0xSI+ZcBEYtF9J5/6egrEYuAq2oWRQRJX11QH7PVLCxcIjur
8Jj2UAFgNVZ9nO4VMry9FUL95K7WfsAfqKBMFRlzC8kPBNVyN/P3FOZuk8DjwEUDhxw7QqtDZLQE
DI3G6hFnMLDDuj4IrtfA9s+iMBDlh8ibT2/42uSjQ2TwVa88fYbIQzsFucz6GHtE0siiinsfGnta
VlgU2A88zoZN1SJqrI05dUDphd7c7DzvxlQuP4vEzvnBvP4b+eUtof/3a2bJh2ID891EoTCwmtY/
I5W0+YDyQi3NUq21qy7+qqiR3omXVeNS8yHLWv9jdmkmBRjHEQ5p5clRN0OkrDM+6vVVfAfqRnai
T9COuxYTwD272+7T1zH66xGk7h45fbGIGwYkp3PrXOXuz5zMKgTcGF6DOSSfvjIjb0eyf+m9aZUB
V/9REFysn5q+GbIeui/n7b+zmnz1CimB2PcfK4oBcq+KgXq0wcIvSElUeB36J7Jae7MTi9WNzotE
6y8JOQsOAjg4Fm5vbn+bsRWaBsR8BZYzjyRT/l6TEXHvEE6xUrSoDmIyPuk4sZq8PX29mlfR9fIY
Op10jAovwI9ZP9iXWHKYNVWVA6SJlhTW37Oma8ecAUVC1z429VX3s1/EstLgFWFx2EqjQDCTeN8g
W58q3xuqJO2dNsBOObx3sZhfL47djyzn+JzUi18Rw67d/dzzlWqxMV+crSUou7imsnZgYMHYyDCR
1sI3KAom4n3JjY9EET92Umtggas1kQXwfWd87/gK6zk9Yg34BfVYd6pFaUvTDSushU22SVrwv5j4
2A6dabambUIYRapxyk0kPWplkiK2RJRyorT0kYcJa7KSiBj+m2tfPlWUT2SeUpabBrFTxwfA8pIj
7Q6hdexjMZao9nx8wGWJvU8cg55SwsttubXrMNt5NveJeE0Br3SCz9fMm6xarYIPYX6Uez5udSx6
hegY7vDAD2CzkUHfKo+/wI/P8xTFayhFwb9B45QAXNZCIEa35oiB8QShz/rooQ0D+RDEHiLJ1euS
mSNRosYpqLhYkskLN9nEyfbiu7yMHlv3DPZdI9plySEVdywOk470obi+d2BIuDVV8SJK+Z76HAX8
2tLwMKAZEsF3DNR2eqFJ7pt7e3PxfNCIzA13Qpu4vnNCkpswJGJSCoQhd136xdnLbMaYjveWUlOM
4IJQMYyp2mL6uoo7iXwTOHbID2rLveyCFdyfpnj+jiX+42m6ZAqQb3DQWOhQjBAtkZY2WstxaZKX
n7+1a0UPfdqpIoOOM4X8IsPtKbrE1TRDeol/mPqII6TToyiFk3RUAzH8r3OXiJD6Fsrb1ZtTk+hq
uuk7MtYz94D4sAuljq/gOqgP3ubKLVRQbXI2QEhRIcSJicrfLj67wDJLpfOh4PrDUHtjiMFDEZY4
pXE+6A/E98YEjG1E7wl+usGQBWep7/9uqnWxZ08v4Ebowe8TrVm+yAR0g46nk6XcpHZcR4cXF1DK
h15sR7VO4pjgBiJnS6K/FzmiWJWfsq7310hqfmbJ3SApnupLH9uNQJub/uUAlF5QPimH71yg/ctQ
mCL1b27mb0s2kUcR3bcjKLvB3Qhcp0/AHysSzpNY0QsI+yIIwIOwQLttGo4H1a+/SdtMZLmJFXjv
ee0rC1lhngljGQxeDKVEPLHzoD6kmCQrgeWtTKR3744wEk9+ENJ6zboe02o792pqM1hpKNhiX4Po
SDtrKBlhQEZErkEUqZMuYuVBpSPCFoxAPUJommiHfTtifYrjwEhcZ8MZCQ9EKj25PtahicXKy8SW
zboI+rmor0k1F3MdwsyqsZAin0V9CrTjab6XeZzav/YEEmK97gjo29gKXoqom28cXHhLS5HK+RhW
bGzqekCi53Ad4qC0c5IqlG7vZGw63w3XNi6ecKtSPoXSb72n7FXF1U+yfpVNnubYQ+BRkr3DHN/b
tBHKrRjElhsrzui36Y0uxv9uv+Y20v0mwANVN3hWRBPoKCcFYNfOTPzq5nhI8lYC6lRmAsOtoI7T
5GK45iNvI7XTVEAFg8aW2+mpTmvSjzMWjnkxIacmlqtzjawlpf/qV7i0FQaJbf1mLOcurqwnG9QB
9nEDMHewVE+R1/1VnvA4AKBwTPTV6TgJdi7/m2xSmGRt6+Dpni8gSS75SMpVHyTQXe3PM9EhBoK7
HguFmCntonW7yV0GLF8qXi2Xkofw571ZxIOv+qHAjzdobS39FG1JZthYsvY23LrWI+8dHrYelUJo
2ZHtYi0epoDGinFSg4qVWFP3MBOxyw64YwPcwTBmUDCg4hapcQQEi+u8mX3+XfDcX0BNSgifNFOD
aNW1sBLcBr0qsblBbUso4jlR3gy/T1dAhrEY1Gw4U4KPkyrF30/U9zcUV9R11Abu9BLhBqoRztbK
mtwmDlsu5zH6deqHcFyCbEIR1O+UZXV9VlMKxUSkP1gLkwcvtyhaQTrga9il6wkf2TizswZkayOs
LTDLYD5guTEkvPX9KU2SJq9F9LF5yDNa6GtChfMuQEzvxdjUCfOawMCROvKM/c2XPmvGQ69XU6zc
9KUlai+7m41UYSqFgeo9Kyn3ofeNT+T1l1c6BPOKhKiODkv4HYw8DYr2sSj2YwjEyvWvkR6RLgnE
dFxGsFPbL77aCheX4f1oRk7B/F2ttmMskIicbWkWoAVS1NTG4MwailEictKpSw2UB0gIYkSSbJdj
mjKnHR0cEK4XlLvpX9X0HRseAMmhuo8CYFhYzQZwnMhgIgzNXMZr1IxidCrlVlSQ2OlW5SrT1dQF
x2uUT8Y0O/Mg/9A3mCpeeteFZrgGwe1yZ/oGTwqwP3ytXg6fKWS5WfNsJY6RTDfahw0X3a23PLFG
fiq+2GTPns+tI8O7RRj1u6djfTeWiUWtQ5zoO2/poHUZmRZEXKgb3Hze4uS7hXuk/uPhwEWgNRlP
u5B4YDFY23HYCMFLHQq4uDiewvHmlaqmYzWnbGAm5h+pI+tEaTdo4I3wKEJW2SxrW3bpITpT3HV6
xe05YFvnHPQAcBdpeRR93bP3mctBAy8D9jBxu4uxUWjXQ3IJw/O3hNUkqaPQYpdw9a1FRpEVQp02
a/qXzr/Q26+T34CfVXElBn+TC6HVzUsDmm78VrlaxGq17htC1uw9QV0R8rqRKumZ1rjETZXeZw1z
jN+cAIUsHsUgDT4voUy5xGRYJAsikWgfa1YUkxElv+n7knvbAok2qglCa8/+DkpU1AvqIlwTagFc
hADLQ5HFFCmUDF/s5OMKp/b9qvl9nngZ6VlnH7tESakMHUeQmwhpK9aMxw8JJJeQknRVcZx0PFyL
oBQ6Zb6F7QbBHB6IYO2Yz2BttT/ahMeNUUGnr53U7FVBe8oGfyrMkf5ndBfFZnF5gLEScZXS19fj
oRP/rjRNj4xl9fJyB/V8FgdNylkmPlpBaXvtfBqM/zNM9LLU9d41aaNu+mFNq7raFYW1dHnRlfqx
wDswt/DL3PVRA0rrj2hXwLso5hy8YfW9gX34WmPG8gtPr7BMQV5pEUjQ6W2Pch+gUV7weXWFSsO1
ViZsbo56UbwAirMbmIldyIrCtVB4pYqQFlL50xUlhc6NI3uc0LWxn7JZ60vxZ/cq0NKHOaYmYhXI
2ghL0J1/cgCOEPPp2kQbrFTQNxvZRHPlL/azv1For2GBjqYidK2AhXG0FSeMUfLEEwDswJd7ffo/
abkLyhEL7pisOJKti0ugXJQ9/tvLK7jqXZZAUoPSnlNlMgMRCR8jew/XfvGc7fhzhFDvw5BY3hpX
j/dTbnUVkNrHMWODFW/qA8kHiufxVh+xULm0cds/Es9OZEz7c/1Aby6s6u6S6iEVeVuf+wKYQWTL
bTREBqpA5danK1ekyK1UIHSC9XGTafA0k3SqWdVJg26NFfM4UpclZ1MDsoDJVD7LkZZlk+oQsPJj
8GKvNSXFY6tnpbbi3AfKFgc0bqhRrHw0cuxxjmHiFbxd+PEwJdWM5tXyXpAC43I/OY05Ceba9qeW
6u0CulmwmTU6vx+E1IlgHCQPgN+6eUjNCwRBVPvfdHhYnnByLF/mUDpeFCLRLrzpwB+FWhj15v3v
LTL8+9NyzKkFn3EhXmqNYiR7qbsJ3R4+iHnn2rpji9ppEZNuYgGTXbh+9LMP2zAbJpHRaoGKavoa
vU0G8vQBFTRH8FX7/sV6EN/oMehCixxfLCrtQBQR5Zn34TDsxxblUt6yoDli5PkCWxulJ42TRaRs
hHR4r6cJ4ZKrGETRtelriNVaurhW923r+THLCqogeNq2PiS2BVCC+PAMQvdnFGj4CvAL0/+ZuCiD
HRsRSmsmoTYPbJYRuxXtN35VfPoeePGs09mt9mh1Te/d1dvzyr4mLfNS+MK8t3LZYrGs3kRwbwNb
ezPxfKhtTUfWV5lsWRt2RAP8iC8OSjHF/B4TZ58Gu+a/HECBRCjEXPnl8uaPIGF5Ha2SAo0/kcUK
hdTCnqqJt8YKmzEEnonlcwDP3ptgjZIO8SBCFVWI/fPKea4XbQFYrPDrlkGsqj4RHBy+/A4VwVqm
iHr49puvy7IkU4ZXdCrJspLOHxHmmx4rnygrom2pIMWFxXb+q6RSjShgh6argEt8w9R5gCpGsMh+
XIrsjBmDy2aIvmaH1JtkaJGltQn0LKaRqG0gF2bJLbKs9t8FmesEpsHxG7AV5FwJSa2HbQXKr0Pc
W5PpCBMqrBcbIUZb/EvrRA4wBR92f+L4HPv4Fe1DvN37mAHz4KCmen2m7BIJodhp5fWsvTCiJ4FA
mVxTz4tg24JtxjH0EIAZGoEy30XzYwwkBlVrjB81aDSwwHUuNJzmnYQ2H2PfbXY6qDMigsJMKHdK
h+c9R6QXYnASeL3cVzXCBw6rtpPhIBKryivs1y1naQKAFECxu73fQpnYiFBukIDiCF4H6zckAttM
sP19Flk1zd6sFrhKv1nH9sEFT65vCThJd0wJArnuBA3BtsBeiDu8TRmk10iBRZkIo4/uBhsFS9md
Q7J1NoH/92udhL53caTIokjFb44kE/Fy0+afwSDqTbzWJjaCICcUMoHYSF1aBP4TLKHOaLfKa41Q
5MORxtajN49k5IMqIJA1K6ZEI5u3EPsiTkyk8MhaZsOJR1l0yPAwBL1ZNVB1ERdy/tn+27xoyO1l
yiezxZ12eT873oY6bxHgeUdj1qrvjF0OhQw3VKpQ/50YoVFZ6VxgR044unyckkWI3n7iShrKiOmA
7SBBevMuo4vORYJt4/bv4ylwwGSbd1f6E9H9dYjFTW9g85bf7en/6kqmqgw01jFpIoXrU92BG3VP
6U3jP7W2SF9iOU/Lt/+I+oD+2helR4XsKvt6M8ot63y10et19vrJcDvlyf1nF3IUfFv75NB/t9We
x3JkQtSzFm9D0ftgkup2DP8dNP+PigFhTMzOV8gomRn3vSNtDHiwwr6r4rsSrGOAZtIzt8QXuY6p
Xm0/KpGbC181bRlVO/IbnznqvPmJ7yfGK4I7H6mz+bcCJPPwc+RdHHJawMpj1NDkO7Gvu4+mXGu2
/ZJQr4ZLEeC3NPpTSkBJklTD3DMyGOBVWU39e9Jwqe8IdHHPJWa5GD3NgqYC8Ak1XQu9WH/5uLtb
XnjUwi5BnYxUTAo6E2iWKU5cekgV4WLJsUabQyArFJhbIwo4zJz6ysLqO/4MDPi9QdHvr1fnDbtH
zvZLDPBLGFWGviRidyWgOGbIM3V/SPs7fF1cogjLI1iAfd+6LlBJKbv8ft6tmRla4maHUbf68PIu
3rxBwhNCNhypV2o9FyNtRxfGc9yYggqRJSy+81Df2LKC3TCwmm54ZNfxHti4+tH27zzysbGUeh+0
zJy5V/YtAE6EzJuQ5XJirXsOU9qQ5F4DBeR7yNF8f61w2aq790rgYBm00+ASzj3AUdhIzis7rnAX
jDUSfNKttL+VzHTTpyAn77X4kcq8TEmyTt+i0bkrJD9Ao7JSDE8tHMNLpr5KbUBkQgC8x0bA5Xox
LuG0j1+YOJMQgf5KDGjm2emmtSxlvaN/LUZm6he4D8MZtMtAix2pJF5jyTt5vrGCFNYj15qPHEaQ
m/HeAHMCgb7U5Eyi0Tc9bBG/+plGh8AdaTuxsz1Qm4ljV5lbhOa/dA7o6piMpY3i4O24Vir8O4xB
MnkqqeIa37j/xn6VTEofr5Ie28F932iTKdJbVTu1xpRAV51+RNqCKmGycPxDerL0vx/eOSbTRvqx
F/4r+WVhGRj5Xzx6pwkRamQLTLFZzSKE1e/D0pGXY44Sp1UaYyUZiwxImMAfgWpafPDVrL3TRjOm
MNn3BJzW/mTcVaoiWT3yLrRanJKAzV036TvEl/+m/Jv/OxFqvEaAg/AegKWgRMlvfizH4zpEgRTF
jq/BZNQP5o2Ha5Tra6Nfa8g3FxgNKMsDRJsE8jniNENzsR04cael7bmShnu1UbSJ2JGHQy9NGTIa
xprN3lXM/y4v8+GlQ83nfyCxj4rNplX1cz/jv4IIAYGkxeERJ/An0CiUY/gyzJUnpu0SRvVUIku+
1aW074C4U3Y9YSHTBQu+wkUbHyjy9aIH8/jjUklvdnS3thTpHquFuNyIYTEHIz7/S/pUe9Uz+4Uw
n1meepoRf0t0A8+KOAC9vYC5oS585RWNDm8Sx94hzf/YvCx1n3ovwJfsFB3g7jmdAjRSWYy2A20u
BwETX+Dr7HwYPOnbOk+uz2Cj4yVz+0/dxIYKcXWy0EX6/+ur5pbHdHq/4owK38cx6zkd9102DoZo
MgBMOSEm9RlgRGGoqllRfP0s+ZpRnNf3Cq6jGHoWuxT9y+I853nOPabFdamPSkCfp43a7+Jc3ftM
VmThbHBQNt2t/ekN/ghiOcqMkbaNXf8YmY+PrXh+HuqjzA2jSoXMlD/LLT0Urz7ZIq9+1XU1otUm
7ErWIATudxIaWGDhScpEq927oQnnVJmXIb7C/8eyOghOXlPTjKWsZucc2hr/HIYCDb/D2fX8GsFT
LrZeTHRsjGTO1Cp1MviBRUfrz+so9qrYADXt72xTFI12uO/bcTqf7VoDP0qzuu/9VIkmmwDxOmgs
P5cjWxXgAGx+dXmScRdbWYRD5Q1dTC1USMYIrUIRYRpUfkWr5D4sHO+eInm63mrLghJz7D4Qgp4j
xbf25yOqnyv3Xirg1FxvMhzNynAqI29pL3HPWicrgmGU5hHJnOAbjMJS5DFrgxtShooThQS8ezHL
NF5aPPuh48d2eVgSD1a8ItyBmEfWXErwIbzaGcpbb2UmwqDPaobwMQcq4TWJqTesUpsD0P5SZ4JD
t8/JTnD2Tv1zczywYhlJV0V38asK8cZPCa56Yy7yxi5pCJal4JSNk22JCCiCttcIB0DIbxFkGZYG
xMyeV9A2ehQn9M26V/T+1vhnusdYWUzrMUonHIR0HsT6Xjhk2Sxupym3hO4y0OBdhKsB8CEW9iVE
1Gss38yz5E8z6QiXDe/xm5ydTIxmF86Jtc/voVQpv3XDjvC2cAOwT+VcDnynPHgnl8oeNdNWwYYV
/SZ6GUIeOrbZuHE36S6gbGgPKWezNTY86Xd2vqLpIDal3SrloU0O/Lx0k7VvsirUhyoTh++gd1Tp
Fe14LgvpXxD0WFYCTlytpZ1Sm5CBSu95RMOqpO7baFvWUmJi4lug8fXLse6VPuIyRMEot6be9Edz
UBaNbOlMqjqOCsnTgqiJqHwC1VXI2tKfaVcBYDid/raW/uB/eh0t4vn2HYP3W1M1idiYYvC2o6Ma
QVmWJShWCtuPWYiauKecrDLDjwXSwai3rjMxGOXMFEZfYqW8/0AQ2CClL8iBzA1+iva3YDJ1Egkg
QwmgKYU/brgedkLhlsrN6FDYD1v0HaY31Sx4Z7wzXFf6Ck8eDpBFV+B8HqwH9tkOj6Io35+bnGNx
dgzqckrgl0h4+G1fSexZHpoIFQ5RX9+QTyl7FwHB2xWdLE1/7UYsR02WkdOEg1fjhlB79yzlDouf
BdlsKzN5FoPz/nJ7poKDey9LPvLcbhD/WlEAkYjrjOdm2SbqZ4s8guQvPcgcbld2HOAj65bvApX2
tA6j5N4yGexWVewX7/2r6R+RdlFJjVN+b2rF8nkQRPpAeTvtIokzU+0yvNUvuPIeno62stKnXU5U
iBr48VQjoLOEmnqItE4hpfRXHMGyY2uGVB4jVEkerDkYrVXEclMLN6aRx+s0mKaIv2cWqPjAO98q
82RyyGcYWbXqYTduMmR2L7GDxKgWIQiwFG7eexnyrOX8JZVuHLU+X+ambi/cS4rjifxMq67wuXUe
iwjJBlSt8YrfI8uhgjXqXGj4Uw3Cnm6qPdBAqXPb9wz0B6jGlB4mauTAPwea+Ckg89mISSIaUeRd
U3nwLMlgmr7boz3Sh815lsVvz8FIiOnk7Wsy+FfMCTAnsZcVlXFsFEOAbEav/e4Cwm1Pp/FOCP5G
paK+GOSoy7hhqpaIv2LRT2PQTmbU8qL2U/EWIda0Sfi7TGUXoEirMUxBRw8Fobb5nbHh22qJ0Q5k
oUVzEGXDjRIoN3C7Rni7ZVwJPmaTQducZUnRQy4lnsmM+N8PB0dw57nrLjp7aaI1QDiXcgwgYGHl
9WBttEWCzLQUso7eJTATQL3gPpUa0SZILUzeX1j54uYhQybRYntinSkIDZrfPuoQdjiZ41/YY0ME
nmBWW3qCZcXdZbtsPF5EY60CZr4TiFBgtQvXrb1BbW2Hk6q0+WJRKiNMJWpuTrET01KGDKhEmN4K
Q1FqVxMQjE0CdMMRo2ErfMUU1Smf42c7uki0hO4zLTMbpm/dDE9/O/iZE5/xH9teOTasjT/Vmb6n
L9sra8pfXt5ZcOqMj0qp71bgrneQJ4qCkBdc4TvRgRF+eH/FB1373E+X0vjEscrbVV+7rrGL+8JY
fzULC+Im39NdxIvRcrdObzfJyjcfqsn2Jnl7zUeEr9Y2oh9I8Y0W+4ZJyTaFj41ZiWuFeVdM34GP
PHXVWx25nH/nL7vs5+whhxqyJxg4y/bUqrlPH7b2YZgVJeIEE4d8p9ltSedLIXCij/WC0ulXrEtx
p7OkBoJvfsDc6GZVdNSpAfiKJliDb/AF8DbZbE7+y0UjjWXs/8CcLm+MyxcnT1dhjqTAw8EcsJK6
Tb+nKm1P5gziCcoDl7vEpNvvP64TRw9bbuexQ1t69tOO53DKAPBSCLBdRwtHNGyqNAaXh0YJbeRc
PVHUJ7ULpDK0DNYwhd1rs3yJbhbH+6u/zZ78pn3zp/2XBYs+R49LrWl4f/Q8Ixg7pRyIBgJv+hNU
Mes2y0ez4uIbi+Yog9E+kzU2ERQH6+WTLyjb2tiY7PXxDXe9UWHlitOEmCqFarJqbwo1rh19/ZN9
s0E1rhHP87QMj9Yo9AjluW0EWsecpa0GWMzT1w3ZqEDalwqmqZv7hP9RxmKLyBszoEzY5aKrQv3b
NUUqLLJ86EuHgA5gfb4hsbkJRA7U8DJThPjShgsyQy0G0ER3ZwNgfhg/8BeeyDbhSUSZQvHzOuO/
M6JqWz6FKazHChKx6mJJofQ9WFDfvG6rFdRoIhZcOztlWtxM1aTlD6DnXG9MtiPjaSE2XJxCmWXT
B1UqgBWyrtnU7pGa1uMbHrWcmOwZt1xlqPPdhHbuiaLiwoeao6jorLqc5nWyAcEcyUCJdJ15RS67
+QsokD4xr60SLJr7BhlCdzQ03ONslZj555GOleHFM6MykyiNxpbXzsUdf0CGfzc9uHwh2JTu15Yy
qXZwcOpxUgunYsIxXn424vn11Gxwo9QsvMmOg1hsAngKWVk/N2uZqxQbbZUqWIpLJy47cixiZYAr
3Hq2CdFur3xn+jgcDpSiRFPMBJzkJD4ytgXCmpG3jfLIxY65rlczLMudFOA2WUsFacrdfVxE4dhQ
fDB7zOgLTcphHSIn5E3p/e1FbTbHCcVlzcapKU5GU/pjsnJGmzUoa6dZ6gJWe3ukfJuh99qa5/ge
wY+e7Wkf4BdfbH8BOpacQNGQTtYOL29+7e0ulSjA9BqKlJIJEuooqayLmhCyoM25GhGLf8ukzpm2
YgYHC/ExJM3THbar9FPuJHPlwV7v2ozDhcRsSUpXJmqErAsX3CGMo3vc5x3hm2CYeEez/qdMpXWZ
U4S1j3AYJW11TkyfQX+ZbE2Y4QTdz8ARhbER+/LyLDrx78ssHbd8x7WPVDw71MjLILpWFb+1ApaH
yAykV8IzOpIWNgXywt8TPHAXq9GMXseuG7mfVX5TK5j9HEo3AYac4JfvDiC5Ayw9U3F7G9wsVXT8
jDjn9x94frgi+Br0/u+VXOoMPCo01fIbytpmGy2G5R084qX0FNZabqeEQyieFhmm5EN13L/SDvgt
GYBcnXVSFnuFApuXNogwkieTDJMPMVR/O3fONY/+UjJRkyIaa6FVEyg9bCJHo8INP1fk0q26V9aT
zBPUch4Pm/X9n+RiqQBzPGsH+QRycdFylLEyHfiw+9cFX9EyvSe1BpiXDm+aFt59HXRzpZG9OwsK
U1jNfnAj3XbeALZMWZN17SMlHvDmEphrrBxXlUptZq92fW3ZVl3+vUWrUcy4FAiY2auMZLkq+9pG
pOowKqJFJQtKdAiKEKiNQycGzw/rhtlraxB1ncLRd1BsVggQ5dTM1UIZgXTY4A5XeopYwemfPqnx
QhrjBHNeggUl/gaHq3jsOx2/CfYdlWtSpyIz/JuU3UAGxJLzsUBlCTOa7ywuG5nVYO7lKBJZ+8Ft
8mmE1yACq4X2+y9NbB0bi5I0exnxuUHCVm4RKTtk7tcQQ7UoHv66vOVwFxcFj7uicUEYe5Je3Lc/
A9jpY7JxgJBgrqGlQb/ealZKTbFKqNi3MYzOXyMP7McWN/dCTonmJdt15ne+98I5Zp5RCppGABPN
CXnIV+D7KeS9zJwMKy2VN4wEEf91ZZmFWsGODPpP++INfWFi/RITUx1UYD2HIRpklLlMxeVY3CpO
sI9/R2tVni+sC8RVA/SCPn9TTd4mjOqAv1Onl+gWU9JwTqyPBca0nt9klb6ZOrGCZ23L0VYlcTLe
vlWLcTrX2+chaVs/HW1q6ckOEHRPpbMoreyjtVFY685DHQ2M1cz69vIp3LOLX1bGcnEjNZkEJTIN
4j2qIjztxr66eMbVfSTykeWkdOVz2U8lH6/ibVOGbxbUqvIreBbdalN0kH3r1Ks+3LWNnsOh8aO/
VK7rUI9T+uzAEciPY6cS1kgfjDtWuIKbbLt95H8ZXUGzZcECBuseaxbymWtuziIbyqaP2GSJ+r+y
fgVXSQUqlQk/t5+cLT7Mn5ApL5SQ6OEyvRgQ4tbuJmTEw7AD6PFUqlExU4UlnCRzym6Y6rs80Ji1
oIp22N9zjUSdLsBigKZi26Wiix6DTsyrguxbtTaCOjb9bYVJ31IH9hXo7Oxo0zV5t/OrWob5qwhD
po0XlQmcoDqvWrWWtO/7ANsOiifVd6d2MkoyeNoo/X53sxp/ONe683HCrjSUqvvyLOLIEHvcX3fK
+IoILPfPw2X5PdcWzm4JFPcM3e7We45GoCfpqTrT/Cl++XmzzQj77slN1lYcdNZBsJUiIPPeVei4
iV5s6OcTzpgfhVrlZX9rwbOVw7FQPvsggbmzpQh3hBpNH4oLLfpQfxb+GQ+rFHdB7TwqvEAmdPVe
zbZhESHZexVyJmkXtIvOvZmcH9A/TgyBRUiHWvr1hTndzBrntGj8RN6ulVQSwslOnxSo5nKx/Oim
XIpLZ0Kx4E8fAH1R9NsuKQjcfciMYCeJIIDvEOz/D03QII9paaYXDAEhHg2oJD1JGRPwSldAWrsM
bTYNJl5HK8IP0DUwBjyyFQcBppPfImfptyg2/PytvntZDjLgcUcjsEu0I2mOTt7oPnrV7WdsI1Py
ZODbVemnO6rlT1IBYZJyTN/AAm5k0l1mKBCcdSzWzjZiGKP8eJ0r++TRXbFG6bsQofx4B6c8m+Nh
TbTh4QtVpxdeIK6PfxTdaXhQs5dDMEj7FtYACKocOQTYvOV3D1TpiiTk+kQoaoFU2KlKHoUnq6Yo
btxiVdlhVVapLpuHK7wL0WquMoABT35znjSzFsLpdBgqKBdRpDfkxkYFBdxvcTVPAMs0aXB9zbM3
MQr1rmluoGTTe400ykq4BW6a3ZFwfsRtwy+280YibkjbRyc2nQPvM3DhpmD0dKvjRjFBZ6F1z5oo
vvAbCemjUpISNdxbxNLs9dXV5lWY5ETHdN7cw/xFdPWxXcu9BBcCdM6a6ip4T1Zikzyx/doqyF5t
ZIo2W1kPCd3+7RPgD+stb+lez23VOE4/vEEgsaITZtfXRAtJyZEcSLaqdDROY31xjlhBpd9mNUln
SaNYvWIKoiesZ/QItJYOUdRh9UgoTx+FUkDyKZWwQlWAFR6UU+gL3ncoKRNrMj1R5Gj/Vd/rzWlR
o1hNVsch78rCgUPBdWCKls8NOYGfwvUG1/evgrjuR8Q/CPn8VO1XD8c21N2o1R6L4LfrcJf3Tymm
m9CHgb02V20tHW4Rjlxq0IWuoU9fD4cKkc036ii2zGgbouxEsjSOVE4aHV0CmrSR6lwisNK6loiK
DrRNa6REpo6x3Zq6hCxEwwF/2Ikor9Q1DZItqN6XO8gqEEflf336XOdna/EbwozX29YKIGc4xwI6
7EeWS7AFHgGpr/iYpiSaFN62UKey637BzHEFbAsj2Rk9sHne209Ekq0UaluYzjSaB+wfjeQKxqZh
0xOLylpbTWplVd0SRZXvzawV3Ij4ei0nZcPm5tNzEiiuaXwLVXVnMl5UwcPfr3zMZBnZDeVpngIa
oPY/tAAWUa36gM1cq8AASxgBdO5B4pEZeUih4RZ+9o8s6y6ZtAADWTJgdWItnTj6L9xd8vUWiGp2
hw6egOHS7yn643REiFNrSMfdAszaxCvStAG7rnUljWyUHWk+rOEtHjO5g3S5b5MRgtQFTH6T5Q7x
uvw4nwssylQFR+joix5XtddE+VhfQ5FaRVFNHLgry6klBD1tq6azDtoLaOXXWcVK9e+hqTm0q7Gt
dpEI22oeRDjtgUqgOEkN+MgdioRLjF4QXjt4qtJ/qA98L5x43yz8xlPmFwhUltbvky0d+jwuX3HJ
A3esnpJpoGHQgOI19AxXE9p9qvC7bzGmXgGi8/R31ITZ1j4nfCF7YRiGIvg3Q9JEOObUmWq9XI0J
7P6uOAbv0fEKd7p7VXRX1p0ZwSRh+/kSndPtUhLxLwOiP0Jie4VTcgFfLW0o9zbf45+Q8tdv1/y9
kCdO1NeDDKcJ7b2Yaq4hAkxwf9FcghqTfsmPoi1kRqeTU3ibtW4vKhIcT20uigq1+cBOB213mhPF
HAYrugncrBtYXp9cWsTee1H6KJa+wjk96B3FSfHvyFoxSkZ+1Mwdh9oY5gCQSJYwlf2L4HwJAigH
4eKcQFWp6R4rib/td1oSS+FQlDiL8J4DlBYqJDzRyNArKywdZPSdyUYs8r8ZcTVxSlFGpGlGl6G1
qMBunSBGHo6reauOpXL3D52TZlhhsf+tsINdsB0l6D5zM+fBOi8A+oc2+tMPk5YvssveYdDxqB4E
2ec86vpkKo2kPoZSPWAwRl8sUec7CiCsNirbkGc9YAdw5b1Zics1hhT4HDYGhaO7LLj3qTRcBPkK
5/XZ9Cz+rKSvdvyBciT0M73tvn7S41uHLVW9Ai65ASvuqftQOEhofO0ajC6EhlJDOLrrDaW8zH5h
161x7/9z5uf4476U/W6Oz+x/d2xISGC+oqnqskR2H+u6ZoyiAL8joQJ2t2ELcO6+brkClvm4bUax
a7ABhruR4Z19iys93W9qWsE1PhZ+gdvBVHUFbTkJr88W3tnHO1se2nwfuTBOTV6OIldnEPm3F7Fb
Rkx0GQ6iydykF8XQzl358mxqbMY4MLSYAAAlZcJsyG4/3Kea+im+BVglYVvLIA+sEZj16rMQbDTe
Halr4fDQ9/tFHLnaC+aDPjMq9CTC/dO0S/hoS4GMRqYyTiBd/gn52ztcLb1Q9hobqcwBI+EO7V55
ebJmQo7Fja17wbKThOhvu/7KMIxEkNjqd0Ek0ocOVxYMmoB28n8+IKMjtj5s37gCANpsCmYMF7Yf
lGrd5/dHX7+5X31Fuaemgd2Z71Lia61CnClUDtOXqao/mud84FmU+G4pz2c50o8uBgUYatcppSJT
+3bVeL+WTNoKY9njTZpA7h2L0Q16mVE56VED21wuEhO4PQ8mczOp0t4MeNAJ70+6XtVhY7fbCcsR
04UTP735J12BwEPaKPGQ/v5cHAd6QQ6EA9LR/9vFd2zb2hL3WUoI8XTSXVKM66yx9ZO0n60zacji
m861uaynPMqvfJ2oow0roiICmrOYJDfsJI/QZ8kY06FUl5nLIX6XBvFtVnFTHG2+tUQ9T7RSKwwf
vJprO06Inw9aZQVaNx02Ig+W88AsamBfeSi+AcGNuUVBeKqsMV0t4hLzW41nqL1JIpk5EvxwPT25
d7u5iD0Af9977dwADJ6lW4XuCXuhbjyUZmI5ZWPfWDmwUKLu0zOGAxHICtKY2f1GTkk7qmrKK+ns
NZfkAYARpinqNgOUx9UMyUKBuqkP2Mj+BwImx9kssdt6hqmHWT74dAQ738WvhKTxUIaJ026JVVmx
rqXfrF20ZUzdE4AYNMFPsF2ry8FkwR0i93gj3/lI0ubhwu+JSpEKZPkYI3jh41Md1cT3bh0BtNKJ
SUTp7lo/emeP+RSONoVgivKeMot3l9HYmG2WTBo33zE/AoukgeMq/aMZpvd/lQ2TbjVOVMltDUIw
9HqtLmwD0ALf3NRMYv3dAyzblhirUAchmD4pEnwCULD6UZLBuVAuxfiJguJ0gRF7Kug8WbsYBd2O
uh5N6Lr0N1CW9uEnuRGl6VsYQPA9eUn2ys/Fz1T7gfcprMisLKzdS5nZ7u1Coc5EUXkbagksd62f
aczvaxFsZ7DNXn3Utd82FIA6lvG8ZR25tXCs3InH2IIHRFb6FK7RZ5illPpRbmELgsJsTCew1ibV
7PI6eQnBwK8eGWGZHs7mE6xtuu/7+rI7KkSxzIzFa0hWJTC70G+yI2yuh0MIqHnLYK6jR6uEciQj
IywQhv/cdMeNi8Et89xcchI6ptDUMeVhdH+Z0v9T1nRCSuOg1OVr+NNK7Vk7s093/9amXO3VaIuI
HbLV4fGd2tqEGdKuja65/RQZlsOa3o0eEinlrkIIW/zjF4SkPjZXI14CZMXdHTU7Oa9ljepG8TgX
CrNgXwtRKR654ox1S/epwKvIeGTx9pMJ1mFf5nYqKjVJWqgWbBYt43byHCQdf0z8XzNCUoh/D31u
+xNAAAkRCSt2k/HmZd8KNeLZZ1YRKvTZvwQ87OkKKCSJTKsFTs5kMtI5M+r3hO7z69ovy6ouWgWk
It9xEgWcQh7ZceMVfSnVATQnW/k6MoZ7p6odQ0bZoubBFnuS4pVGJDRmykcvvNnRBh66H/V96ec1
scxVUkB9/q4DgRPyMT86OfeRpj4I3AkfZH7x1KmO7xBeALeBGKnEHOS+uWwiX0DJa973J2WTkvj9
E8EvfTZ1d5nD+y+WgnYdZn1dr5TMJ5vHhdR9Pj0TjadyC4ME56WgG3Wv0JC0pR553N4qzZl8idFz
/U/eN36OPId+vtJ1lwjz+z0uAItrfHn9vrDll7eIYwluwxXyuz3n1oj5muaXWjdmUe9zm0URl5qg
aFlo5ECnl6sMkyu87wjBK0U/2Fkux4vCjBpD0E34jhfFwOlsyrcOs0Q/LjZ7v5zdVKOSgFMP38F8
T90xjvuJtChb39lQ3yjVV6sHr8ePM5b+GX8aWBQCRb9NFt0CATs7AIyJDOUMv37q0aQ/cD4J2+SY
GmNqtmxNvEoVIQMwpdy5EeQman47DuaC/P5ZDprF7Y39KewYb2viWRIgvkMrNFtzXt+x9NZKgVkL
6Tvxx3rGIOSj4Lhbf7CG6hz0caOhxoANC3E/f1NMYEtxbZ502ZmBGsh+uGrEvff6K8Bwia9+tC6p
o5avNfccHoQBj+i5wQo2em/IFbNz4zQi4jV3TObWluB+BgdAD0Ga0DTwjieXjSyfTbvIIuQo5WQS
INEmU0azltUfDmfOA1S1GhTMqHZnUk9M7SgnYTqHJGV35hAibeE6jhA8UDkuRU/zLNRDsmbDl94a
4kcmckvxehniMN3L1zVWCIVFOWGfFdPxzklu90vHPkzUBjZOg9wo0bjHBgqmoZ5y1KMI/bFyzzCS
KvfiQuw9HDMNt1NRWpD5YlfbrvSa/kfF5LwrpIpWV5jbACIbalCRD9J4EoEBmIMGQ3AFhYOMNz+V
1euw1Go/2potFX+i83HFGsVeihmaCdYlyZGa3jJnEb0EUPnlYMq+rmPlVcXt9IbZJMgEsDMK9jva
JqOvaxMMi1LDkvRcnkdBjNKfsocBzNrrJpVDAXDW2tzz8HJdd2aHN7FuYdsDlBTqbBouhVw/Pk2X
Owsa9H/5FZNfFudXyG4bNW+edsjSijm9J4AAeZoyMcItIqSuHxjjbAJ/kxdNEdzyAIoleFRedmxy
JGFn9g2xL6a7YW4H6hmfkB0Q+OSF58esdtsNLfcUyAbcxQqwRBMb17gpr4uGqzMmw2venYOKwmzK
pDtdBc6mL5NQ/Td9Jq/RGr/yQL2Tzt6X2aM/b/4Ulspyhcn8XCkyayJnGHdNwPNqcfRxMwf17Mzp
hNbukn5zTT3M2P9xeEJRXmTUz76b5pDJnm+qQgFT3dy1TZJ8uOemre/DWXJ8ZvXNwAI7G2PEM8cC
TBnrZVRDzpm2rrMIs9KS16scIoxJT/vWXMKAwSmuTEcQ86rLBytmmu81ywKrcTUkh0Ckj7vYCHUF
6421bpsf4hSZ1vbHumbqkv33DJiuo49LtTpPBt4/yfUgVsWyfy8JS9IAlBpGvSLJNsaJ4uXwcQ0t
U2B48JZgpx0UEFqCz/4LJcd4DD/1cuh/9ACI6AkbZZKHrj9U5CmOUGlQhSvpbdmDqt+QeVwdvSBK
YsuXv8aNh8SYq8EUoVZHX51J6YHJva9e1Tm2EKyggmiVfqbDrWVHJDWiAc4frPTGIJm5jP4bxybw
hGVZHcyy46I0Ci10YwyEMhoz7j5wpCu5i65X1ExEiCkV9jF7NErve5u9a0x+CERIqq2aRxj9Wkwu
vURcL2DnWC4JvlN+q7mgNL6YG0fiS24+h+yrE95CYHJgzh0e/+mD6mH0gqwmTot9jgm1ZhLdYsF3
bCPwUN8daTnFdZD9RfuadQKkfbhaVj98d3XwFI5k+pMJxnSEkwHPQ9LBWkpBw/sYArnQhkLc1R2b
i4gE3qo0Oj1OSEgiH6aaTqK63SX4zm4H539to/GRhiCR/ZxnkyoXtIoSV8S6pfb83OjIG+oVY6hy
ZQf5OIEjZUMEAvjGHpV6aod9FFNDUZC2CpVj4mPq8e5zmvfGvH0oApkTaQQuXQXif9oeMh1gF6N1
tHA4vJEEMr2ffKDBwtDsULZfqOT7hb0G12d8o4JJTRI94Z5nwTFCAuS3h3i/WM0UeVweEv2yzLpD
NETsiWBhwHIG437X+tVkN07YpyXt8nNu5Lim3dAgF6JRATymVku+pAlDIbrw94nNN8psr0eWosyi
2oEMSMzSUr9PlZ7G1+Nnl5EBsWmYm6x2gc3TRcx8ScycTxpfZWeMNULH4xJXf2/jZjPBul9KT9Ow
wnCzAa07EHleTvLSaGec9/UNG8OFRbNDgruJZgFeEaBAPhvZqLlTtEuyRKH18G0oTSZYYm4Sw49u
AXKeH74bR8ZQ/rcL54h/DeHpX/AEKfwvmxf5JVvExtCcctWceX3E+N4gSbjbMEabSHhDj8WTMFxb
ycJddm85YY/EL8amEK7ABEJ9wva275HzWljlGvkdJQfczH3xwoLm0a3gGJJ6yNI7xobE5a3JpoB6
9t9wbAjLIgo0T7fWRqfqoH3iw6J5LF3srplsCtKHKiSEXHes/ulU3ELNsz1BJyUg0HMB8F/6X+Vz
Vvy7hW3XtxGZKXApEvNIMGCQmT/++vAStKUj7LCtkHXcxX0mUVBQsxNj1LfyupNDPrYBdtNwL0aL
AumtzGVO5c6+dXnAMJt3j4gAmrhd8Ovz476DaMRzxUIj93oxUMNw+hcOYiz66SVEqLOykSLW76ff
XE5OkdLBEPJbmk+yBQoOb8sB6KcT0oGnUxdv+ZaKx8HbfR95T3twEUSxhvm24OOq2V9stab9j6/L
+AzZTXS8L5S3Em4OhyTAPPKFaHJuq2QLgLnyNgHdEqktZ57anZ3n7YCYH/9FI72/D42yKqQlOpkg
j5muWXKHm1FTpknapgroE2qlJaMGzvRmwn5l9CweHuIQ2VggmFG8gw1elhSwWhjC4ptLfUvqvKOf
VctBe15dzmP66I21RvIwIqH+fer4stWn1yLnOU2EeYj7Z8aU09VLY0eVHdlNPCIGIJ94NWsnYOVv
ZYc44GpkWl7gePWwzLxWHY48r1epajWbi889wKAbN521ljnAv+pkPzFps2armHd80cJhno998dIO
bgwC5UZ/JR8VzfmC4oY30AuxcSkrRqCQ5oYFPWXJx0pSWBX8lG4T7ltk3XSzgCS+OHwEhIo7h1HC
HMazMyjXq01sb1kZ2eqFG516HpqXTkxsU16ZC4l3xIco2BHbAzXsyZLuZ7xFHZWlYKVDhGZja4wn
Qp6TpOwkpiyXZ2n3YqZiUmCtEOnJ03dfaX6qQLrzDZF2J3YB6ay4xS6hIa8kvSmtWSN7ejfMFSg+
/jZVXPZhEUMJyVmWadeEuDXwQjzA1BOFF617RSFNf8b25UDXHROX7m89+ZYrHg3rBRJvtHMVK/tV
ufxBd8OmVyt3+S5cBUk8wNdsFxsbSPm7K/xNe6UlfG4UijF1L5jI1S3umH2lAQKq51nNBMGE9B9d
kPDYyyRYPRPf1HvGiQg+YVf28VhlFeWtnUH10zAFNsnDERm/OBaHFjCfcbIrQzm1bmZspDiH0MAb
2Yr5y+aS0kB/S1w5t4u1QxWDkyymLOjKVSNpB8yC4X6FXXhvq5mHG+l85EVDd887pb+La4Ed1ACI
ddrKrlcKbh/ilo/kCJImuLDm3ZDMUu6dJyhtGv+qIiGMTy0cSel8dPoLzejFqoejF0rcL5lTMOib
pA2rgMO61RIgEN8G/bKpiDFpp5H4tvVN/tMsD4/Am/7nuiPuHenCbrS80mC2YDja+tKXkS5GY8Rr
h8qHsw3DY8B67aj6EMxMsxFgMNVLIZOxSa2VdwlIGvh6Z7pVxFgKbPUz4Xw94aqMAvtPSuoi1TY3
HSS9p+bswO4AMCFIWOlsAfjjBcbByU0NI2SG2g1ou/l2/ywTOhwbv+vWVIb/jmKyPnj1Z+s456Fp
PenRrqt7EpsvqcbvBO07JKqrV96mxMPB4MF1JOz9BJXzgJuxFY4zPWKRgHu8J2bmIeM7pTzUiOLG
6FxOt1x+lGrkmEVuHI0O9u/qcij6OzcRzffkYGFrIbJ1a/ETJwxWGTG8HzNdHEcXkddPSe5H/cti
e9kkvF6HDdFzK4Oy8JYuLnn3IG92WH4i2kSKpEnyJrLHJs9dTJVMP8sBSCwANidSI0J7dEx3s+fG
Kmxm18RKZ8Qf7+2nlp5Dl1AsYnMS6Suc+dfI6XQWaefCVoDMhs0b3N/WTn00IuFXtHXZXxOHYcWN
BXFRA+1Mp/jJmKt0KqMoB2x3t62FwmiU3UUz9kteyA9DqCoa+QUDtVHjnlMRz42Euv+zm5VFUbtG
r3JtgCFE0WH1sdsoXdsuAG8R4vnC6li33pZR/YYmp+mBxbz+nMkCFhqQQNy8v7kXF1rW9YHNDTG5
IdxKw7nuNi6HsdAw4DzfJ/mAn//cx6JclsUG8MNs0qCcrbSSqOBILLRIcmJCSDz+Yx8QG7Z91M5X
KqEqNvR1k4R3Fsbxm3fD0wLzikZBIuydvGDZiKZhmrOoerQYZHHksm9KKKH1s6RSU48MmUOPQVi+
kgzJHKJC9zjut9SGy5duVcI2A7XfdjOzPcq1YkbQsko1sxXH8akhkLOHqnxKC29uHNUByl67dlli
4VxFvRDBMX90RT8xz4R0Z/rptIoHcfJoS+XnqpCG/zLHD8ozkKtQN80EchsstpghBs1IMlKuPPH1
l8ULw/tAj87oUbCfeBxmTWo/oW20AjPNvcylMfkoiIw8gEqgTTJJJV5rpqjq3rX7sZLVrewZhzSY
ePGUIdQhUz76RYQ7yTJLgLwHEFikkglbvS5hJzzbqgdWg6an0HFnE5qQdKqyJHnkTW4/gwo9v6h6
cB9cbWizEgKRd45a5BP9x9v2wYw9lvGaw0FeKIQ+75xdyttNOz0nNZw3Ya/4JhBVwFzMrUg3T1OX
cQiQsAASyz/5NnfadMjsbc+ZAqWqUSfzXE7+cs/2YsJJOP5cAoX7X8Ods0BlNfA7/GXoMTbiK+yb
Z2ArXAvbxPA58ihGCWRBY0IChkHkoMCpcvophPFSu4bs0iB1MKS9kTda8KNeW6EGKDJ6cvDOb0jH
usipLBxYQXeR2MiKO8nOxRPNTl/pIhcizmsAt2iFEp8w01TXFLeEmTvxTgd8v+WSlfRWsYWm7BhY
vpL4utr73WKQ2G3uGhPZEk4ltfEn2iTWp7XC9sWK8PxbUFZaON7fdHjMqie/ueNgud0Niyz5ixMQ
z4w/AxnJnwokDZWNDA4+1zWGpwZc4kjS4GY2c1nJF3XobBK+Rdxqgbg+9aGjBoUjZTYhzigT/L3W
6mbZ3pQGmH22CzsyA7lAqs7QJ1OwCTJEUmwwp8BX+vmSPDODiwITySjtVFGOg4k0+r2UAcKcjwHo
iYy/pLyvazJeplBV/JrzdjNnQvfNRYjn8xxn+b8QD0CO6fF9uo1zzU0unafS0bxy11inAkAxTwSQ
CltZvasVnnOzKBHB/BhY4X2IHCEG+q4gvqmXj7qap9tP3M79JJS7AXADtUsc7M54U9w+Qr1ZSRb7
6lgwFFVq80kkO5LkzKFRRklb3YfT4NrOgTugAv+AztCCQzAHNOuJZLaNShThQlfiqfU79OFFOe9V
KvJLtkSM14TFSc9sP5mexv8l/qzVXwmZdwNQtTUCTX4cnj5oaiUUsH/4nmjx6+VeaB2TteDBTBwJ
Uyu6bI6bi4//TzAcgTuI88T3JYIlyBOwWboT/KecO9YBIDSz/WDrttLEaBUVvfJP4XoKxgaREuON
cXCe9shc0bQT4RzNFKxaPr1qw8rbIOF0y3ogJVEB303pa4wgieolI55Qvri7FF5kMF6fHSwBProV
oXN3A/EgLSDscjwoWvg8NNauFtvs1MOBdyLBHzsWpMjEUXuVt+cxTglShu9AnnB8GUsOlfqY2e4e
JUJMhE4R+14fUSMNoSR/C6DXY2648Wya5wT8b4bvR5gcBH0lV3SdHTVBIhXgjb/WQ9eTCo0ZDBGA
j8HX/uResvbn6xo7zbNbSylnEz9zOt3bXh2/p/uaocJNmF1HQgamx2VxGNowjkRqVn66p8+FK+3+
XjNh/nq9tsaOdxL6cwubyHS+vRnCcWo4927FCxZf4/VkxtKgH73aYCZeNvQ/rn7X/Vfuf2VakAEh
a+dt9CEG3lgnmLJrlG1OguA+mTkd3eZMNYZtTxtnkYsJXZ+uzrwO4JthGJGk6cRPp+F5z20d0Of0
dDikjWP/piH9SsJZnR6LC8n02Bz4xkRU+YsRwn7hbXxcgs0BcZEBe1VQrLBaPihO+Z3jPltBehSc
GXl7b/sizkNqB6yTF0CaiquuL17nTZ8hdw7JdOtrR112Z0FIWo3AEcRKz7fQXvwPZ0Rwy6in5YZt
b94afM/QC8sgmTzKyG0RhV9/7qyMRon+LW8MZLWOxIUMUw+pjQ7rkVEk4J0MH5qmPDYtDnUAb/C4
E0FhUo5shVkiBSJzFla5fzHF4/uPlwLJv0yObjlCHA+b1f8EqUWJYQcE6Bel+yDwvJWmGUXdTvTe
kagbAbSFIm8SbLDx/Fq2KEsUrVhK0lSe8xYZKtFEs+X7nJqkXgfx+WdPceJrW3ATRgt+9eZ/rj+u
5WZN+vuSYGC/VOnNCl3L8e9qNnSnVG8N3wqAllBNWVG/Gi6TKlfbJ/wVkvc45vS1YiCGq07QlyV0
TANu0PZfU3B4emlQ06sYFcWQZLf2C6xpsAstqPLnPLXDS6ysGZFi85KND76DxjgPfXJaPVr+N9oc
C/C3onnbRWhPFaId1IPlBmGdgF1IpsB6iCHg+K1BnSbCrrOGrINcXUMK1iBm65C6d+c32vT2xTnY
eybvn8lDVFCF5kasJVgqUeb5PQ1//6Z+i8e3hmBHtUa/1uNV73/LC3+5QGCf8fz8Ypc+2VMg9u82
dL1GdOFmIiDv9DsmO2lwZBHAgubwarRC4R7oPXWEgrs5org2xRszkojCfaR/L5a2LtinM2YcQ6tK
/i0qiiwJSLY7doMH9OmPf6LUafRxp9viTuErxk1cCvK7JDY4Ndu1fGz6AXj24sbfjz+FadSetPyV
qxIXyehlAWeanHBC3qmY7BGz8UrKlqf/abFMdp4ff+Myl09tV9CzvPkGH9wfq86YG+2wHY5iMqJZ
y+49jGbn3T+ztOZoTn03TfwCDFpkC1khQUyHHWchnx7s2unQ2j9a+ZsSrLfTdqpx+N5khHNqbTFm
m9MDgKPpiUXlLgLhd57suurHq7/4YrGpvT65qj6HnhF+/2d2DUNRqqA69rE/yd9HBeMeODV1gCWX
esCtTL4r8GvGFalKZ4ViYSszM6/fCOY+INi7R8TtGgtVyiF/iWhg71oX/ws7CEYPS3J3/Gb8apUS
dHm23iq/uWSLGIHIaXMzcDYB1vXFY+uO0p55QEGOJLHKKE+ljaW1JA71dsnxuB0EX5V9OqYKgB+v
+hxoVXtCCA0ogFYm8gFkpP6QuQlzgici16zvxT0XW/RDEDnHuPq3/LA+GdYcSfBASlgakZ6ZFPM0
YlUqNXDkZAisIUWPqUGnAigt+ZP8SmZvT5iO7zQBUxGBY+GE8wlefm5pUk0xXg7me/bWdkfvQVZg
r+V5aeI8RGdlII965HOx+H9u/yYmcBWTQPQsprKAn3+Hw6bFUfBmsdAsWSI+pPuMWy5nfGuz+hpm
iXMB/FxjKDN8qyG3lHeYMe+yPUto5F+RpGfEwPqXR6q/sTcwlF5+ihuYjPk9ZWIowpes0n1reSdy
5sP2maJTao+05ZZYEfxH1WV8MnA0gaRn5qDJSSkhjlNiuHlcQQmpN3jYVGtFVPV2PjUNfYay1Tfq
KVIfYfWge9e51UDin4BTzB21N9aWp//NevZSIP6ODcT9RR29IWeOLge5PqxYxjVUhTbbFjfVHGJm
NsUbyPhY3CEngq3ywSLFUtr4pXxUCntktrMH5qxN2YKzDsyBr/CNqiFvei9LoOfIgptscRRgyp4X
1Y+lmJhy50P+Y24hZLpwxkRli7bN8gLA1RfTF5fm0M1QH1mbI35mON8ceu8ULw+IGH81zCXf0F5q
t7fiTEr20Y06sZrPlITmcgi9TLVldhaSKk9TqmySip5Bn4joOvHde502fceAGoIa6TcG26ZR3GgE
c1T16cMdtoLsWU0boaEv+Zjvjry8OlY/r5zmhOd4CeA0wfHW9vvfN0M+6fARqY0a6OCND21LH3Ig
U9eEJipcCgMhLdlY1xtnaqe/bhCs9CiXWNll5oN4F4CzrKCE8ZhTX9eKz5arp7dsUOZlKiORsRyO
uCWT5C4dM43Ea4bXHT1Hop/wD/7UUEQE5CNjzuzhfVENYi7738TnqcNep/JXvQWXlMfSOtwfXKut
Yr4t+ArE1eX56XcgWN1JYQ7ERMydKygasOw+sohyUBQ2qE4sKXJo11xNZlI/a/7O2r5KUaka7Kq7
MpWKlFyXOeURquZ2zDIeCO4P8Z6yOa2jqFyMkUut4BRVz9/XWpjuk5GKKIvvaMahMYdEk0JehKR5
wE7VblRJbrihkM19wRqebZGVdH/fAHLkMP/FzF7peaZqBQ1rnDuEQPdppt3QH0dihWsGZCRpWvL2
UMFSt9ulBm/NEomuJI9FPD+R/iklq9z0NyuLMWjU66D/o4keyU7s+Xg5OoObY3ORmT9XnymLjMnB
GD+GT80dTxq91tVSFVKOpc7PybuD9pvspposefazOJLN3V4sn8pAt5dbpPejvBxQQGS/WMoJ45iQ
Mfu1GX6iZyor4pUB589BPBr1shv7ykpKMyrzaWVnGMRvaUCNYgLFYZU3+YyQgCmiMoszKHXwNKZ4
9clpmKfYS5oFT5qg+AT6p6m/K458UGjAXEmzLgNl608X7lX5hErr+1p1YsaL/ZxXRhi/HsYwuU6O
rTWLUhrPfyLEgEH/3tyhm5XomW8r+p7o+qeCQU4f/2fwLKxEvbg2CvJXiXavMCZCzXdWXEy6t0lB
Wm+IC4ICphtgPBUegsfVdsONtTrwibw73/8YN/wMI+AYl2NSpxpYashpG8MTGNztb+Uglxlji2i5
5gl85a2C30gyhfTD/DHkCRxjvuzr4P5VgYAnjeIrjIozN2Y/b2MAjvAcfVuIIw8bH8bVBBhRLkD5
9IdBPMj9ti+B7wuzFiBKrkAzVXD3nyjX/rw7usKdwLBjmyaJoDS+XY9E00MbukwrkfvS1wO7OQN1
Nsum8YiL00nvRi2DrYl+6zrJk2UkwzjrcB5jZWk0aRyf1QjUgnbOqqzoM4jwuZiwU/+HVSaRM/Aq
o9iRxBP9vKHtPPOdyfo6K/p8KnvU3jkyGFgMGya+f7VnrG6e5lfClauzQPbAsGl3r5P25ZdegicS
VpQbZyCPRphqzGpzhkBgrwhUDITxEDxu/y270bP2SNZ9BPF80i/1CvQ88t3YOOAo5qx5bun55Rzl
li6GuyOM9qI9XTTXKlF9LVj2dYWTMhLx1lVP2+6WNkCuB97prowzBtlyGIbN/pwcnBVOjoOQTcTf
8SS7MauWzCrBuRV+mHCglHMyhhuhsjlZ64vmmQlDttMA3ybLvwYPekmrbBcAvJQBu0uxInVdsKPk
UQsmSbjMgDMjQ7bMiGys5vpRbJfJ3SHnf4QEwX/vPW418bfsJbWwOrzlW6hmNQsHGLh7oCNZI6Qu
H70mWkkCnGxEPyYGta0e7I9wTolWbr7j09KTjtn4h1H27OcQ9jS5UFEV5e26yQlCM9cnRX7mAbRl
NmFIqiwUKtCSXupN3fgSr2OX3nOXt1sCp2amu5GWUD0oDFMMenCtX2tsXpybZ+qLH4cWvAiP13Gv
VBK2R4HIdfTXQ7Yum1W7aHpgv0SQG783FHqw74EipR38zCt0z1qPACHm0kwWCiuPL30B1+WIMDZf
T6TwF7xbfM4D0vQYNpamzrdcsMf7ScsbDnaGItxK6i7dQNQIlH49tzF8mgnylmx3GgYNXIJq+Xpl
mL6iz6Ae0mlqmddJgkUAL0rjJ5A9TxTefZo2DJeiXgysF25i9rx69FwfQGOX6TH+/XU608z0h2e5
e2j6kefsz5Pl7YmsoITGFXBofJEsvT0GqVOy9qCy+3oL5uGoFR+3omlUOuaLCm/xFxsc+XVlplHO
zeUC0yBHZ3fvUfswwXe7jF9YcBlG07ZJH3VQ4rJBCaNAa3TDWPBJAAvUIIIq8XAp7IXvuHMJFKN4
tcniNzB24sVWvpR3wCL/Q8S7BBOt6DOZo6mzAJ9pSYU7cUE8FvmNbyb94Er3Ys9VI2EWGN+qpF+W
ZxtqjqOriU50rshPBRFvYRjZoTdujOJ4/gyiKXVKnPbD2lFtzzplGveROEPTHVCUgzrm9XzCIzOB
GphX54mGE4IJpFIjwraB1eUveNhvgvSV8bLRWk1JoXFMh0j1Czcg638MceqCtwBMYeb7xkiCOcsw
m6+aERXYkjsJo2nVxpOcTECVp+jCdD3/6EPe4vUXNZ7sGbdjQEpMb8a8553MPYWHur0uB9BWXSYO
LicbGsYknxlmydSVfHaTHE9fgOXCx8fU1tIGSGigo7kopiaMoeUMKWmgprIXzP9Du0R1fqY2lTZw
np/zhtO+7KM1cG8zPBlH9DMdF8xz/SdUaLHSwrTxXycOtV5DA/PSQE8YjsPm5d552RF5hdc9bcEF
FDTrqoGv6ehrWwjg3RLHjrLoEA0FdUNcECQ8duOE0yA5jtapZ7uK4HQo0rDH+5Up7QptmqoeZ8ZW
Ch3dzCrHNMa3OIobgGEcS82bacBCa2eQFsRkcjr0SJMz0hzF9p8jEiJN9ilum149mcrGkGcM6NT9
xBbTpoErZ2LSi7lLfcN6dNW28XhYlb2Gskw8k9fvOW5BXP4/rfp/HINHIyjS4giLpBXi9xgM0CAK
bRnjU9nUKf2EyPK1I9e4mhKPndwQgv8XIYq8eauSY5VY/d/YMxIU9GZToI9HNxo3RI/+8v9+OSu+
JoYIa1mTaARQwQ507o59/ryB3JdmZOGs0GMdwkZGnpzaWzw3m54f0GzND0TcJOWwQxwvSSReIWU9
D17yguZEy6Kn2mOsNXM4kjOhxIhWj54Sdptu4nGfkmDihd2+hrwHhM+t1xiLh75XzwvifQTsEGX4
YlzIR7HNYCiylGVHHkeQC5oVEM66DJ2XYEtRr6LeFP2NWSz0ZPYw2rOTT8Seii7/eJe8wLgjXRID
tH82z6ZVk4gmcBiLWvBR7AwqJ0aHALWsWCfPSZnv50AXpNbJ4AkEeRKiGnNCp7jbvMBlCfVQiEl2
P3122u/miZGY4jUcESIgSqZLE+SBISdxEERY+tlK7Qq76/O038LtFjKL0XcqiaoksJRm5plxmZnf
GSFYZ4PJSHliUVG9eQVdxyxlDU9e0RKzT/Cu8ZMAt5lx3EsOWNUIo5/CiHJVLAAo1btpn4i5avEi
e/vxbPPFY/004uvyxfm9buSqZz0LO1nFBwTLdY7Mulnnhe0KuGaYwNKQgfbGU7SPSLGA8hQ22R6K
Hx2J/r7NQcuW09TkF1gwbNQk3YiHesqbU07kPaVwqcmBgy1YcPiBLuy0QQpICZ/k8j/Rvo3wPINu
1cF2kU8QHDQkkmWSBGq1acm4hA+GMKlyR18LpLGrKE4ILpdSnSQ8XeIWdFEJ3whOyjHHi/TENkDA
r/LdEhjtbfj1Ja/mULcprhnmNXXYzxp1/rLSZ7wROQIdQGAQD6JzPcCh/GPYB/DR5z9E7+O1cwaY
0EjVQsTDNzNR5GeemTh+p04z6OwcpLx0/5x6jdw87FU8fPIQXSJfCE6/OSOPUv6pyCuZO34l1NQ8
cnqJyCo8VwLYRGW2kFx7isfYVInuM4sN3G14L6sIpNcfVQheJGM9I7RncQvB/R50PUjJTYaEPtaq
G2PcuUxh/KB2WqwPn5XdofQY5RoVDAsYp3yMZkkHWY0hSbZcyZ2/R6vhN8u05ZNbXVsUw4sT/v80
EuV+JTK7DlrAqAAf7LCR3zkw4R8geCqhffdGetDfNu6mzKksabVIG8DSCyac8a5ktKRjsytRWBJF
evoHZ2InhLSvB2X+2Jn5HQRxr9QcW7umbtIh+Q4nlZYDQvTl2FprpH1oXAtHXxHjG8x4J8BCjqum
C0IfPX6++TzcHwFFycNlNg9n+NqEteuLdt9+4k7gsrjXpDPmzTmADV4FNEV1gijs4NkgqlWqvNMY
HDNWYm029jsYLSVJW0gUBz9oOjwda0+cmbPvhqRKKvoTN8mQSz1SbUosRS2JqSzLmXo/5Dx4zcon
Q8EgN8312Gnw98pHSHxXhDivIMKccjmFOqXCJP9IbewkEGw3obBuah9M5A8zSg0q316EbUgFFVS3
3FnS7hRbDU1Q3BWLFbnYsidvLWJ6IXk7LTB75EaDbw2/bqyXTJKrpt28QEiaoCXUYm0Qsfr0oWix
CpL2zSEsri5PaGoOd9NQEDOhLrsQdbbcpz8lUzJZNrcOyWCdYRvzON7ZPN+xJ028O+HwMpSLoHja
rAOZlo7YMBg4o7SsVIsm7n82cobCBRrDZazreVzF1HaNOuNcKJ/WRMd7FjipGiNw1X4zC9K2CpR0
t1PaPjQ6Lq4phej3vGTZLOaeR+md8YOACmMpgDu3c5BaMKZREpRJVYIQaJ1XOPwrXlJVGaRWiXfI
ryY2Q5C9P+ceixjlFCEF9rZ4w+GzPV6+gj2czSU0z5jelMlnfcacfzwD8aNkiH6ODDAihOmDqE7H
gOeOCfYqDSkvcKtRtnD0RVjmoCbxnEBFzv9xsWROwLPvtFNHfLScYI1SOGgqkTyeIOqY/z7rSmd1
FDZ9roY4b4FFWXO2OaQYDdHE3WJzmK3Z7tMSjXUZqMQRzTNeI7KkIBVWpgar0HImYezCjRrp0wP0
L+BkbSG8qgBALz3sYVG5q/L5X0enctS304aoKLdSWgzWIBGDQON5dL6bxKr04BmKDH+yDF4coBbQ
j6IFIobIILMLbw7WRBMED9rHqSfNmQwwZ3g0dzU9lD9xFhzV8MqVd9lw9a713GRn6MQ7ETKmE0au
l3+EKbnrDlcoJHO4+5NwTjnK7d+imoizOb3sXe12nIgDXCiJuwXtI8wwwgJXgTdb2NNfsV7J+L0J
hITO4XCNib/aR5V1i91i+edvKkocbx3EQh3XzTnvwfUR48usJxMh9GzBY7cM1azNpXz8TGvEV98q
ktqery5hHeAFjE/6xD3jiKtZC+Nm+SQhG4KeKhpnEBY+PN9xQLydMblRxdfGjs3m9AR4oifZun/y
dNqI7yapVeogfpn5/n0+JiE+Z9rVcdOhL5j9W6iYdKkHZiQjmBDRtBUhZre69Hfp1io8pzxlEXXB
ZSExRCLpHx3YYAUh6iYpT01sVg9E4hOV+h5kr5cd3euXwdUc3ZdWA99dCWS0SAcD1XMMomtd2NDq
kMOxDiJQZULp5OMaWwtZp1/7MQ1dpGJB4AFIUvW/gl8eFCgqXyIpHAEe3Wx3p1d/yxy+vBrcvhEP
xGjSIC648BEMeHZ/Vo0ws/7MpUwQIINP3oIp/NpAQXmoJPvo0KmcgeBtU2jqb6DODQ42QPJ190ns
lRMU+MZxn+wzQ2c+7nrdChVnMXKHSOWgUaa4nk1AOmx+WbUI0rlK7qXu5cHIUWU4sGPT2rToDxQF
ieNVnJd0g5pQQYkAMgvp2ddHLylwBdCg1FB+EZcDm0y6/aXLuhM7/PzYnhB7F+hLcU60h9EEKnCF
se6N+jI4il5dhylqpo/CQFogqoSmhkpBxMrGpKNVbtrnR2oNrCb+TergTEOMEGMRAaAlbd/8t0RR
oT9Y0I7d5juHLurJRLMOYVwJ2tP+mioa0EZdI6y5EYy4m1ECnbwf9QhgZs9B1pbEB8og+LtmlghV
KHVBIHE1V2sTOw0ZfxXCLFdAGEQc7AaXjAE2lvYcx7/PbLhSsl5oTgRDD7QRSaA7/rHCSsa5extS
rv/CWFAWiV8Vz8Vg8PxUGfqf+0rlK1+fn+IwrrxfXvwhWA+GREwjhCese/R74QhPBlSShKoMFvXO
nK39vyTmqtZM8MD4jE/Em9hepPWu2/UJwp21HWzqGbcyIxnqtE7dL20ZAdRBSbNxnbRBjq4uS+Kk
/w8OcsMWvu/p30aVqgxI9GmHsrE1JoHrpgwrdryWsuZI08PrPtckRZZ577NIImnKFA5jlnLBH7WG
oz4x+aD61Y/kYkVpCcO15LiIxEM/yW+UTphhFrKmiU2hGRUJJIgZzuPyBYgJC1hF11kpq1fQGWan
4ZZVpB7qtIhqoUc48kKaQW9CQR1DSmZu2u//RTTU/fj8PQ2K6ljQHWuOCRjL2KaMwv805EQKrMqz
29ddpFJh5xQ1dk1iu3ge+cPrhrMOZeZ+mWCeK8aKbAr4mzWCxCAxXL6u3bRmYEA6/ec1ZDviqm1V
SsfT9oHUfdB2M37C9BzxxzzYBF/5+DjaiufytIVPaYJIhlDwfrcW2kNbJHu8Ub1Hy6BBX76RHm8X
V1K8Rj0PvG3lpckWKNfqh7ak/EWABOj9/msRQfH4uKYLLIaBRMP1DguDG/BMs95+N5febrP6FOMD
0XGVk9wzIsF5lWjGvRiN6CErBdtjutjWPC6R/5E7wZt489yOGjipUlZ+G0tUVkG88vQVjvywTXPU
ehwzYkLJ42WZD+m4Kr8/XU+64YR+H9FSx8OQXFNfzBDxqnso5rk1boC9EcZR83BYWb7fcRL4sxPH
oht/SXfAnqxfIPcuQCbuhdGQztrYEUgIqvJrERtBzoS4NVXnDNXl5WI8Akge5olQ545mu6SDl2Ee
qZqChdmfcf8hiQCZBhJh/lZUkU1muanE8TKerG4YqCDZpZPLMybwoUSoeQfAG8ryAAroWc2P5ycT
pYAHR7ki3nRv+h0q9Dtm7HMI8tjgG18HKQNyk2WCOhuo1mhRRQX010TqH/90mWGCNTnNy6+hIcCO
lEq94prNpkEAImuMzty0QHekUbZtdOSA9OCOpNnp3T6dXGCOXXn1bEd8uLYzOXU30aZAfcI2Gi83
4hfg4VvuY+kmTRTIeaDK4zYHZMYbncPE1UnwFcw01jIntCw3nqPUmyqDYLrTfympq/NUIPZgR9Qb
u7kYLorh4/8DIpC0oEVO8Ncb4S9XZRD5axVlgLyvQGWFw7RAOrhTpOvrUMkNldKsDetoKTIy20lS
aV3Bg95wA+hy6rN0NOU69ai96nRgAIERJ7VxDXcKl4jp3mVKGxI3hfN9Pn5dfaVVMyE2tvuFm9a+
PAKmqLndXr5eoPEj1JZa1W8YLyMfzobZQvJwwDkzbp2W1gt2UQTG++GiWLFULB0/LAKPIh4epWY+
+sTPArCB2Q28c+QlMk/yMcHbTc4pnhzKeiv5EGG150BRfb7Ram4HRPPUXr3cjVazqbY9Pnnr0pQM
6Fou/kLguXiBe3k+h9o8NZMDhlejgQHtSF2YSumBTA8iOmPGSN8W9GMT2c7x5TLs0mGFqfmWyxrj
weLa7yiN151RJYoJvczbEpl31eUjE5aq04L808ygu8BjKZq5LhFPBjTi2k9cW43fW5W8zWn4VEYd
dNV0wL5eNLW7EGagiv+vBRUpX6C+YpUTCDk6skonxzj/gAJ0BPeBJa+2C0ldV5b37hYRJcVWvXFB
F9iKuW7cMut55kw1mp983G9FeM5CL8shhPZ8M7JERQy5DjbUGLHghNpFYnqBW2VsLSdfmvXKlJKQ
hCe6FrqY0Q12+ExfJKXL/Jz7TFTj9cBh2sUkWpyQYbRgJ0i3y3vEm/TWaIap09xoEu5P4ycHxPBX
PN7Ttta4Znyatr2hP82HT7wa1pEuJrH0TzS6nFOW4fKkvPyzIOOQMZ3MGZoXIIZCbq84j6CrvXxM
WFmpnl5Zg1pOBYRSslyU8QRHsux8Bd0TSRnsjulGDfvKKi04K8BFyLAu364Fl2gfYIRPmJ24LJ8K
4IYpc8JSotjX+2UbRfmoBdTPsbLrSzngTHSAsOEplLH9dKSDNnNnSHk7f+8fUjoKl1t/fEFB3/72
LaPeJ3wVNs4Hm5BCC/IOgIpwMYHi7M4hr28p4GLMdTKXeO9ZlQD5WgWga1uoSAVv7rW1uCyb2QQC
5wGMDGBG/350sjw6J85xf7Jv4iCq+jgxfnUrblt5n5VWxrHT6TR3CdJS725TBcQm+pOi5xNqdSOW
jYoO6C1TW/1wcPLSwgv0ODAE07Zq27Y7/sK8s7jq5p1XlVJKy4FAVrXAnKv7bLkYJ3gd/Ifo/xDG
NzgBbv1zPqkIUmjbVykO5ovOoQPtX3C/9T8GvmspzkaSJ2ptRQKK6+O2ogKdLVuYN62f279xVpPN
bP/MYjt7PFTS2066pAE/j9Eh8xPMsdIFg3ikyg3JtFkMX9WMTOp9PQFMO5+gUsy7hGQHkvMRcS9D
WiOzIm8fr5YXW9FJiK8mIy04eSoDX7HHEyeGCGvSw2scu0OsDlQSTowt9+lHIsxiJw7ZGdbNWiSE
yRBIzqSq2HZXEj36f7NL7KafKbcPovBWiWRmiDtW+jDcg6YLmGf5Tj0MC+7GaKlTZS/SEe4c9AYM
R/WY2B48rXm+P5lfNHCfUsW20g9mp7kOr4LImbVJ63T2xsVnTU/PU2lNdxZRmieudLOO+G5Ioxb3
ao05Ons1PL0oI7XiDui02I87lZqbtxh7TTZlTHlzeJZ8qj6PD2siYkAZDeLFE/avTQxYf9HqFmVc
UEOWORcxDuKLn1vEhnAdIsYGMq4gdsabRZ/eE6345EiLGVjFPlQhxopAX5+U3u1vdH1MFFlFihkI
rtdDKvmouUR6viBhh6khAMOnjFxTMhQ8czlfu7gVTshksYsVzC60AMbHgWgmxsHn721xDLzVxigU
l6xL9EnfmSfnv/G9zz7nhYbrfl1KD3bD2RZnY7GEep9Mr2jRJWSohK6zYQ/OEMaj/uhKsJb3vD0F
RUqnaxPSbQGtqPgmTWk08VsZn4UCfam2/Ir89M7jSd9qNewvUVtqdVeDmzR9Lj7rtLnvZgt+G/VB
wadF/pTmcBP2DZCn+fCZeQ+MzD6vwKsZ/CbvKBzNBaf5zzF6XkmNinqm2u1Zg1RE2UPupbVbszvI
xPyOPHSbEA/HJA3ax0yOVTjcH9sgX5x+dkdJ7zRKTpjomj5x3bEnn27mKms8fSTOG1l9OdnSOsdU
lLg2XITkpJZ1wJF+fDnZMSBdGpUSiXGgO2UayVTCNsXMWG/YSI1ZDd4cu2o6kYb7jmLsjwZagUyP
ERsE0Y099X3GVtzBu3po0p7zhdjTvYWGcN4n3LVJ/xSOUsvzTZFRgA+5vCrq7CHry6JXXR9V5tJo
qFZgy3LhjSjlW/IqR6lZr7cQyCfd2s4kAq8IXAmoBgKigXBHwAK0RQ3KO9PZ4PrXNCsB+gO20ceM
k9Sc0qUwt4y1RolTS+BTyPuFD13VyRebCTonJsWWCou9sViGGT9pYE2p6d7+kJ9zoMRI8htpq0f0
XYLYcUMzms7MAppGZZZ8SgrELpJqbk7lEByMIutZTAY8/SdQxpUBTRIVQe2YTkWrRi3Vni3jdkdt
gDYobbwgejpnHbP8bAWz1L7Zj25Lvn8ivhF6KegN2+BxNPL1zFC91EmeZf+LG/jN9a0ZwV+u1nc9
kkBRjr5vRPmyKvv5KWXDT+he6RW/H1vbZSWfuwvNoWc5ZsQnyEDAUSv2No0V+gVG6Ouzz20ajKY1
IM4DNMWXP9jYlOWEFD7griR1+3wHpb8vuxCnL0ZjsEI8JnImru+5z00sFfRYYyNcJTa1+TLrSN0O
d9jQhzoH1Wwfx5uxJ1db46kgHC9ndfYnQCkqGtrWlkoBkEvNGj9pe96dl/EU7e8S6V9+yZ6ghTME
y5Xq6VxwAAQRTQqClzjf2LcA77TyK/ccPnQb5ZReg61mZB6xugo/IZy6W9K+YE0+TjCLZaxtNznb
VWD/1MYCfzVUG1ZYvj6QSYbOPD1+BBmIbLMOnUV5UwiNeaOCVOPk8zNyOFPXbotXsWyhJpDphRm9
4KcLzsaweh6Okp8jmDthLsBYvbPSXHvpiEyLhdHkXZYhedRlUpd350amDiFbY67j+dVqVg9g6C7R
oPmZJg5Teo5ylI4o5OrQ54CeClJv1vR8e/pDSdPFtuK05T2EijhAWqqcc+0kFQ6QrNaKGh9CC9u8
tgO0zxj47+9rH2tPTpE0/JzKrh07fGuTaKZ+rGw10IT2yR/dlt8zhiifQv7MPJX5uU9ORTm/uU89
G2eX3OUEG9SNHkvGwcw+P7dvJXHiqF6uDm4u9tUVF03Hdw25w8Wrvnrhq/6+WpboRK2m5+HqN57I
UDJ5BGErvhQ8yLin0bcuthgnojvBmL4wzjFh4mLXvcMpeqqLSiBIxIGzqDbA/c3xVeP3PvR3G6hD
Wmo2cU3MniWuLSk4LXI+ugZrTjZk1TaXSb99jwP8eqzA4XTQREVJfUekuJ2ExqKYyhf/JOO3UhDV
X7aimH/dMUk0PBO4PeEzi6rSJ30DdNCiq30ytfsDTITvbs0W3VHVSwbzsRfI5Sibbb1+/74Cx6i7
xc0LaDR3kiMSNnpv63fnKqxP6CPqZ0DM+oe2M8EAkLZThQbiWSmVwR6F69Ve4RipQfrO2TpTU3Rp
zbDGQ2fZCjTu+IeycDaAFQYanmFslbn4atu7NtOqI13ZTtyBYBZbZGJLUvedym4Ek9TwQdkjIXQF
ZccvftKiKRvGCrmVDLn9qltD3Y39jba7vfdDAfVwqbI/C/pUt5DIUvvjT+WhxzAJUCfhx9pmx1Ee
GwstfvKShJ4kg/DNj0t/3ynq8nT8+/7I21rEgcT4vrqvDbGeao/ZSMzPZk6sBfm0RKtboUsMgAO9
lyVbmNZ4VBb5fVMATIau26nXf5xemtkNHkZhzaWyBzCLu4GAEJAO4kqXIKZjns8x576RmuMVaAGu
cDhh5hgN+YmMA6FHCokorgQzZ0sJN88lDVGpCkYOjVGXCKXWo32P0em1orePJjo/zwE5pkDUMpCZ
T4cNDPDh7AnMM2hATAPlGZJ92vNHAGByzouY50tb8FV4SAfy17whVCF2hnVfxyAWZe5Y32nxk/O9
Diaf/r5f6S8BS352au2c/SyLBFDnC15ZqsMpkfZGcYjAeEQwhYKpTCyx8JulcNdsgNHLbU1Fu8r9
VEfEnF9FNVPHPiZO6MT3zkolHqfa0F6QZvlikSIIac8i3LPwPbGg858Bo3RAEiiAR0A46nqUsNM3
Nl+wKxFTze5kZq/eXwJuQShhFYq3vEjeN+mqP2WFwhBJwcts7x5qB/es8uZCdNrw60AOkI//BpE2
4tNTMtGrhxU3uSS7YNzu/z/2cW13f3Ib3Vr4SFCjNVKJiQ+Z00lmB7yTuAxA7bPd3gKxQaNI2rs2
56Ts7fOCkLjwM7YiTEu5zUPBQ/4MdD/7fdt154PiopFZ+hZDx5FmJxZoAtHuhlT+/IDny2B6kqWa
XyE8LvsBxR0V34+/jFQli22lwjiNgTNMlQmCZz1I36+V8Xo1wMJ9z04mZzcZY7LVFFookTOHWSto
VoSdpuUwkIkFYBEJo0rhawVkrohWvNtUqw6KEXrRv8j6sNcs0klYzHxpg5Zky2ym1PQDo2+gCR03
lCn2oVj8k4gXFNC0Oi+clJAslx9heM6g8PjvxcOp0Hkz676Jy8H/uhZJ76eI9kukqESKBXA62iIG
CXUpYPTqL0q9lJVNxdQcmKzwV6m/PvS66LntIlhsGu8MPOnEVnKBq/eCIwwO9fgcBniROvMu7AH5
VwJsnPUO08jQAM+yrTr6o9HAOs9Qft0Lg5xljvRafeeO0makxA7zg/M/STH/MkG6LiEylAPlPhxT
MfU4AiigYupKpj5BG0YBoITBaK43P5Pnm7dkpeHo7pANtaGXFgzlc85+Sij6qYAh7YrgAYup8u75
dZr5CYn5VOTN3eQq1+GfjJFHFL9sW/aG7PMGNORM+u/q7UE98Kl22jqKcnQs/LDKz6qjdf9oDD19
o4l3++eCdkDxqDpbLtv8ekuQokL9zoVTfUFccpZUYIPnhM8RrLkzTt2f5qV1avjo/86omQ4NMWFS
pt20kcwbR1SUmH2o2qYfAId0mWt69oEvRK+zZNH8r1NppGq1et8XEA2tINzJw+2qpSENsoel9Vat
odROe1lBQDVAkwkWoWyzJAslcq2H/T39PaDxABwnXosuh7LjpTOtrITazQM+r5SUhfk2SdWkkqGB
adn3yC9NmfDwhJQ5pu3yWP/EwgcCYcJ85JLtpr5+brC/H48pLZmaEGj9vVVnS9rYMaiej2hvr43x
QZAMAPpkfdjUVeao7GVLnUwcLDzK5PiWjQhDrP1/jtxdmUmBWjuPotczKHQtiDKeelsxWCEnXVns
5B6lKdpYl3mKSZRsFxj5xZlhy58u3b3kyKQ7IoFgHTJDsVCxzR0CggLQzDZ0l38RibzRIUHHZBI3
fN9xMQANuF1T9AUIYQb9GwZD6I4SwVUnUhioXQIBGFt+vdfn1YfL7dNFVHRlvTfF5uxoD6ClvP8o
1pLY7aX2R5ImK2+FwkDmDkADWCM+YOZLuoSIHuNK4iSX83yZswk885cye6WbekGOqZVpHQIoVBXQ
rxr817cds37gB1QOi94T5knUxsDhsoT03TaNCT+UjCIxoT+9cCmJPirYyPq7xEUB3OP927HtjA4a
JtkTjwshCLPS+arjkqWT42WnH1KTVyGQJPdSaiGMaDEHEsvYE/UaMQ66fT5rU8FyXtSCIfT+LV3x
FcirhiPsmUvxiNM7WSVJu4tBSHFlur43d8uOThnmYkivj51durvkwXPBGoZXUJY2BS35FVO/Uuia
6VIOZv+S6HZb+b5amGLIcOxwn4Ey0MPmHNL8dEpOM8xAGkAJC05tujBz2pXcgixuhSaBgMl2IhHS
XZSD3kwMHZyc8pBYKwQvzNOlQeWb1lhgX9JVEt9h4oAjlgUp9CgYu9Ji50QY/THBIAHfEDccz0CF
B3kSPr6ddkdjv2aj+SEkBaIW9XayqYswEAj99/zCizyxGObLYopf/a0zyRT6bohls74iMW+gI7tW
9a8Kv3KwsUv8oe56zfAHCJxFCtIfpCaI79mhYjGBqX71pBVCMPZhtCPLNphWHgcP0wz5BwQmGMZg
8ARFpdqTWtsL9UxPVRm/7WdBwOWTBvZ0/P31933jJJEjbjaCQT+dXSOGTBfUx7rRlJu/dvDpB3yj
rdyN+hyYXgpEFkjOwKdS8Ci8J3SnoJtbFksaA8lTNSVQ/v9tQumRT8bNPZLuFgGc9x20CgIhFJEc
Gjoqweomed88cQODMZ46wzpjxk7QhGG7hqXL/jYTa0n3kA65cwAkmzlyBHmUKKxMVFnWP3mLzJ5D
Rnci7//ZRsTQHnMH3/Bl0b5xbbgQ8wIXzao30i3RQvNw/j3PCkv6XiCRGoGPBrL0Y4/uOr0O3/cZ
GNcTtO8cRt8uBKpxQ1lf1lKzdmRXMiAP0djHQVZSV91uxfSd7ETcAOb97Qf02bQbrtVjCnXQ8z2O
/16NASU8ww5d1ZnOjhqw4w4DHZVFRgj93h7HKp8qAa2RwWk/jzqPS62OidrM1yNY47iYUtl+ejjz
SsVDfp5gNWZ0w65XCsVS7jNGOIAMmPHdgUnDq/8bv54k2tB8wnpqzK9lCgVIHKma/vpdsGOWa/uf
Vnrd5EI50DVpUVadM9KNpiSt3QywleYP1RJLpgRVBD3Lv4QbDKaKNd++4Gl+wp49I858lA6QmZcE
FWbIr6RNDBdrU3GDI7oVCZ3CLZ80/wVcAouhZ+ceuljo9v+GmlpKvQjHHVghV+icgGR4kBlArqSv
TQs9BC/dVsGHQhcNEu4JpiZxmGx+lWdMQ6rFT33jA0ITpUuoKTahjhcLtx12VHCKgwAwp2WKFxj/
meCBnyquyto2j/cqtp/uGJMtllrjMmAIFPq4Q9k8ENyYWz3XRcoOYHGwH4KeQkqSjOzFEDNPD2DH
mfvEunJ9dX03FmTeKzEnyzB9eEdP28l6AthG1z0XGMKPGBj7K60+HSNjfyaMN1cEgfBcl4qtpCTj
JnhYM3D2i0JBPGnIA0IFN3cD2T6DIRhK3Cd010W+/Kzt4eJBHFoJmXtESrqdzyV6S5ASQsdO4YbQ
+FcbrvOKm4IaIhqIaZb7DipxY20xm3qRQm8cZvy4MyldgHcqiAxDF8Z1SfPYyACjfxATn0Ib9qjk
GiIs7e2nlUBY3ya6HaWIpwXLrEFe6FOFeBoba7iJM/Oi8p2YnQiYjfUZlMxvIpAo2quqkkSu/O1s
mztWFq7rNb1yVY+mulyeiby91m29mpU/WJZnnxKYK3pjbQ/+zFLg9/9qjt5Jwrp6Vtr4er4IhYr0
9nYiGebpF7zjLd7MWwEFYvUZ7cJ0LzSqYcVfsQ+YfBrmHYhUjIxc88tqDvzne6rWCqilGu6aXWxh
uWkYJ/3b46mr2v5h720A5TVSu+tvb7ylFHkXRPn12vz2AWYdjbLLf6a26LD1yEwaTkDCXQ8p/ure
Wd6fJid1QsRcqZQjssr6qz8rK315dLYEGmTxu4Jh/ddt9tARER43dv2jly1wbPnBjmw2pr8L6DZN
ts3PMIv82zi9t48BzSSm2tcyneMjqPqg/ecuCe4wwzUsvaAgftszigYORTGOQt9UdOsEx+cRkbr4
UzPy2OKWEzWlfXKDEHKBsZHoElrxJgLbIpBW2EP9q/xKX/gL81qIG5T/mTlOZB3I9jIQoKK1VWQA
u5B5EjmG65B+5EShwVFb/MQ4wC/OYP9Xr9p5Z0NyKl02xRUP04YptVBm1sjGx4xFxiHcZHdmPiTD
WhNGoCvZ+q7NVRTg1mvMteA6u6K87qz1jhhhJtaWFZB2H81dWV+mAkjQxLYrIy1VsPqMcOtVPzaT
OOECdkWQeDvJVOl+V9ngb9Nf77xWb7r+qetCvGcY7LzXWjdywJsnh3LDnkgOGWDr7P8gOPXx2KY1
lpgychfCmWJ8ssbwuYyCiBMTdM04RCdaXqK+QHraRSqSVq3pApaFKgT8ZhBqZXMf6dtjSs6Za69Q
MOYxhumW5TEGlKloismQqqRAlc1Unu5X/lv0mTnkZZhhO5HP7QzX+pVQP4YmuGNsXmsThBTQ0Mdo
z4zfObM2BmIWnPT5askuUwdy/WzZpe3MBMYNiEodB4h0sLxaf2ML7hZvwvpNs/aig2kP+BQK+tFK
jOY5efpDGMN7iphgvHr+VQj5jVTNZG904bN6GFU+GACvJJaDGSn1xm0atDOFVq7ZpnciL+dzG1tj
Q6jKQRR+dNB4tCv6eVHmOadMW3/njnil61JkJDldj2MsQfU4GtqPN1gBUCrlWKpvEJYqQiH3pOjW
bHXePibcicqyqCE+ObL71G5Cx3SOh6cXsNAmkqdq4lhpyM9GMx24z0kiblWnz6k9LM9dbQLPoXdA
yN4vaUYuV828p7jjn2s5XQJKseW4XiwNVpaKELei6YmNVnBF5nANMRcKRftw6A+XO3Bi4g7v4FbO
eMa4hhHXmo/wbgOsRyGURtIV4edmbw5LKPJlothPbDfS5xobBRwjlOC8R+IiGin/Pr7KjwJcqFAi
/3qERoHRYHjbYBEYs6W4lmFzg0hpbt1Yvqt+mGexgyLuZVcyWWIaPgbyCuooaNjddcvX3VlP3rMa
bJRSGpSSiEGgzD7Uj2btmmx54+Bp5cmtvE5O1KBphoNerqWihwhPUBPLS/mcVo9t4KcMYpaQtnbo
Lvhtw4NVUtOciYRJhmgsa7Sft0rgXWhZgC7WPx9UbadNaC49skOf0pnntgy3rjyn6bZ0kNShgf3S
HcIQvfZeyzeDcQTyziDGDQ6OIekYoLZfkbUI942DplYsYcEpmQH3/Jmib501jLpy1VyT5c/oZH/d
Pjxx4WKM86qmcgVk0f37O+S6WD36QhiwJ8HEGY7kvyjkMGe9Em0bHB5TDpjDLQsK8smwWYe0x3Wy
umwFAwZBCIlAsJzsah0S74ZdiN8n0gtaAt1f7MoL0OEDxEYunejr6FBFcKHF4jPDB0HeEhPh8Fj4
ddYZQEZM9flCzIKTSidF9TD7j5Ul1go/f91JcG0ubSqEJiz9FCkemtH6Pe2sjA+kFYWURpmBT8fu
pL4XXgy4ebbFT7ciarw1B7CdJ6NMaAJFB2dOJZ09PKVpbhm8yXLcXU+hSlKRpMc5Cv9KNWp6EVIR
5Wz8S3YDGAAZBoPliUHMBGkiJA4WdFYD7jmgpyOBOFs4TPRcusRCHA11m6HohfmzPNfp7zKqPhYl
8nE3PPyCx2AqympkTCMXbggse2sLWKZbfGB6+0V4k6swYaKTXArDlIUfnn0DEpOoFklGp4dqWUq8
/4Zp2GO0WYdT7IR6MeYfdp68p3lzo1Wj9wdeqGssj0SDOEGtUIESHoCAj3lHBCIBrKQmxrImhvNt
vxR0N/TOxFb7zssdaEb0KrjTHxyNEgRj9MYXFKnsIH6NXACiYxUJpsGdW6MgBgFYkDPt2GlPgSPg
MK0sQXDbdbklUHTuB+I4mEa1bAi70hssbZSvXq+VVsjxFHZ8MDydngwe9nG2rkEh9Rwzc3EBFst/
b0VRpt7iaZwOoE2bv+yn4f3KQDMu+0a31aNUQU81YzzvsetPbxBifKAWzqS6Q+b++OySf8jRK+sC
sssLECfj72/i/ccfPkrnY/C6+n1USVEpsXt67s7uJ3Ro2uDfGsqCTnI1axOL0kWGoB5SiZvKJO76
y49LP9L13bfeenHEinKIaQsVoAqD1J8POxAtqBLIKdpZtGa6mPWigsS6EHNwAKzLkWCshU1ThNJA
un6J/34qFDzAzVZkcJQPQPjIkxTJvW1qkjAiolAXjy/EhLsANzZFR0WgajdC2dgEk1quTApX7DHP
OqyNpaaWAv8N/bZExqcUOEPmNfMcgwbEG7tiavJ3NY2eHwPXtx5cCcsCD2168A92uwGHD/2+Lbul
gLAhCa0trC2Bzi3N1/mngSB6IMlp39QDLleoSgn5NPPjedekO26Tx7qQlAgzyTVeH9AlMFsgAdHK
SxffLP4x8vtT17jaPOSHe+MjJPJZYx1sqMvUbyTIF/A/TSCooq7uOo57kjXNc3u8Qq0fSJxabtSg
QmLXIOGqeKQTBzBpF/LnwYaBdqgFCrwoDPsjCerz89wT8s3ehTcb2SNP4IFNDSVTe6swV2tAOg9X
FyuqVhRvwTtCPl5AAN0hLhDvwF+ekvNElIRERjI6CyHxeuPLOyTRS30g27lIS2tWP1H9Zh6sxHLG
GlhmvATUZcn27W6Tt+YQZl3fOvxlTrnpbCJl3BH7VJ2aj9QNxDrus990MKR3OmztmgeVkpOu6eBn
E8C1vm6QxLRRpcR2ZRwocCo4zFOD5LEqM5gVMjtcdI8pARIhq7sRt092WekVmasCzHv/XgP00KHK
EDG0HEYf6yu3rixdmYcNSjzoydb9Sl/4DZCAJwez+PEPkVWBifbogFY7YeL5okGciT3ig/VU5Upk
AbHTwkjTu5Ts86Heh78iBsfKt5xFM8N1q88b5LIof6sYKD1IA/kBMvT6nKSCCLjEt1Z/lYWxMmAb
LedMntAyL8mD63ETjScFpxic3RGsKn7Rf0ZHWN3jcDlFAKrx1IHn58tlECHJUIcuJjpSYVi0KZ2q
/HqEPN0Cj9PoI1Z8rETfq7vY80fCHR2OQW6DaThcOTDA7bHoqDViZKaSbjCPJAKjAInW6XHP7kXU
SgcOAqnNGOGAcCWge8Mx/bW+jY7v3RHjBCwXNcFED9e+OlJ0kQ9nxh1kGXxoLGCfu45siRlYO8rE
YSC8Qbz5M5optk4Z+ueGfBvnwearNPkVnwjTA/M+Zv5mB1pXvMyLkjVdLUEuLtpoS2A+6ibZjwR9
xbJ0ouXv7s4QxegaVPDFR+cK3IzyxjVsgDAwsMZ5Evj9vTB3qN68JZHqoEwhSegIPSRAtn50kfEu
l1K+HTh0J0ioD8qJPiNLWSTgxqc8jb9LzNsnCujpOwDbz6zxc4LzZTYV/w7HGd+DKt7IK4DP1Vdl
KKSFgfNjRKFr0d9gNCRLykcHUMd0uh+fzxkZT6m5AiBNZEaQlQbHGgRgqPpLbAVZb7oEm5kpE4E9
xBtxMY+qQRv4RXgb6l0sX4DQVTVZL8QmSvbk2u/4mx09FA42Hs0a5nyC8sp0AX+x5MKmXZveIhzG
6EhsU8l5R0JdxA3hIZ/WwT20dykP+RPPXQIfNiomLbqVjrGIG29mS2vqgs0GIpbspPXomu1fA6Pw
TnH8KdSJd7tT/+7f9s8AYBpntjLSewAt8U5/gyJ5FOPDtGNFsYAGY3k4W4CxLRG4/KDReboljO/B
j2YNVbg8qy8DnoPOns2fw7FnJLU8hZ1tUDlt+XvoDunYEsTHJ8ZrUu8DQ/bel+vIVMwEi72mX9dv
r5sGysBMWJIjboOf3wlh3Mm0lWF7xdpQjUfVOOe5mqmKVjYchaeadw0g6VT4WHFMhh0i8OJwJRto
Bxj6z1pWOP7e45tNud/O/Zc5g6y7OCDMkIAiSZm1hIlABanT5DAMNBugRCyMPV4CHABVagvkRXjS
4T1PO5Dp3yX+0cojCEV4+9a/fuJBLXpOta80lj7pgqp4oqLpD2Iz9ehuc8dy7CLXaubJGp8ItsE9
wuAodJNLGq0T7oV8lmrbba8YL42jhT1c5rVncoqS/mtg3deanz8PB6q3xh/UtW2ruDa6y3mRraSY
lBgLCQZlN3pbs7fFNktz5g/gY0uQiwUvEgteLn8+pVSHCkDRfTKM6TGGiJoCVSt/lAEC1htUMKIO
hVM49ZCTtcrUF3NovVieRZfVDf/vkmI2I67l/1ynsKDcCj8Fnnyw7akmMahRzGL04xGcMjBwGucO
r9cZjGJ6PZY+NWfDm7dCFpms8coAOYOYlO9L0Rie+sHIZfwf0JPW96KERwZH4LOK6QRKdn2mXjpH
HHdNlfYLQa4HLCCvWJmSQ11pee7Uqs1YnsEELqsUKhwJk9j0viOL02+YrTSHQF23qmh25reUrHXe
TIW0dH46R+yUvTBqBWVvgIyTljCuJkHZijjIZucjkL3FFGNJq71qWgdkGDIxil8V3KNEXy54tDnA
00Jnm0edzL5RTnN1Z72yb7jsBKpdEtnSDlMMhW07QYSW8hRThWCtdtyTtBUPAvqoWCMmoe/BmyBZ
A77hEgqFuFS/Ji3iNKLsX+j4Fp5oS5GMy20FUiyAcgT/lMA6PaSBx7RCTue8dxvmdLVHE5Kb5ExO
u/64smR7z8jP7PMaY5yQ6eFFppi/uwDGiSnowBP+PrwAflbvkOrga+Y7QsQUgrH+qCVyUlp20iaf
zx3q98EZyZCRqckmWr4W7Zs6+VKz2eidUfsdRLUTOMR2Bz797Sty2HS9A+Gdtxmznytud95zzDcz
S7hN5DQ4oKFtNsjmDqWxqlV/41MxtCQA5SvY/i39ZKuAFhfFQXdFiBKeXxms+AWV66e0x8VqnokI
xlqf66BA/TLSDETI3Ec4kjnRuts7TT7p7/ZVFFBmfRO8HSIo38h0XS1odPGYzBuyqIx48FEn7o8H
+wblNg/h0wAzpJR0GNsOxE6CJzOjR5TUBZEnWe68xYb3GhLRHzRT71BmIPLniGKjTtvZVWKEh9b6
Y9fmXI8EipoHCTQcq9ArufpgO0x8XzdM/hbrKuZb0noHBAnw34PG243Q2AjU3BGIQDDMymqpSIhQ
qI0FNCn6SzSnt2y2uo0wacv9wwYpQY578AmCdP/MWDXJx8wnFs40sffecpc0Q96gGeX06/3imS4E
CobRN5J+hvUcSTdNfGhumGd1HJbOKrAYtLlUNqP/3Jg5yl6s8i/tGVHk+Ch79QzCzi6DaLecMnd5
XQfa9uArKUBQ6k2G/CHqJ+v0UVS8NlhxtHbDs0+/J+SKqvtUPc0NUdIM2PUMDWmPDz853eHg6rC5
00nUiLp3jTv+8quFFWT0cCoVJYCXwd5odJGV9CMCw0GgP1Hb0ABV1Hi72Prb/FOsz1F0eoDsaszo
XIhR/E9ivY7oO04rc8Jp7rztMTRUqc5Jmli2L81iH9/hy94OBVqjEWnHIu6nHz8IUMT8OpDqXMN3
arFh4LPWV24431NAinlr11AL/PYNzbLsr7xF8+EZ4wK9Mh3Ts8fG042IImfZJscLiRhoNCaM2Qcd
Sxc+7ntzwJWvsc5w/bWXqS9Fto2qWKTpZGPWLzn4ORx2696HoBh3ypFTcPj3TxqjTDTrHsqsQR+P
FM05n9qYuh67FzR8IMPwBQOnh4IqybPnzeL63tS1ntQ6iNh7jzaaW3XnIaYV2Qf/vQksNTN7+EJq
SFSmqb2yIo64KithsnOmkhBf4EgECg7hSSwRaI7WvLS7rPgvW3r5lxB75hlgdd0nzOGsdHr34CNC
DlvnTPlmd3IcG08NlILZRsfA/4+iIuXqR0VjY/+UrBGQ5YxD4jhabMoLh4oBqHlTgX9CdZPLH4hP
j+PxV2Y6feAXC+0LFFPvzfVA11BvkZ6dGDc5Fl5fQVwLLwdYz/BTfgUwV+kRq+mMjUNQGWE9Uo+a
NjOCPXRRUIGDiTTvj81zcpayib2IAvS0SdkFCQt+57zmQ2OjjCxl3kzPFz1UeqDcDZIWuY+iad+C
+hgL9LTgtuJDwcioQEH7FNNkzNFLpwLc3An7TY0HhhH+lXrdH7FqKIFIubZg0SXn0OtyeEj/ZxjX
szWnwEuwh7YztCjOPDnKGzKHI0HkynWbAlylx9HdT9IMH8UVEZM2CFmmYBCcNogZ3Eo9a4CRpwc+
9k800YxHD9sBpoVCmdKiyEfG7Xx11zTaJLs8fFqT7OrUBnU7k4gmz0m7fuLXX4VWIXh6vaRtxzSf
guArmIBM7vMs4yKDecQqF2/2MuCcaiqyNLpc6GjSXXWYs6khxGbH4XyOg6ZvPdS6aB55oLJFCR9t
H2KrpNOQie2wFyzWWA0vy8RQmRqiY5fTQ+Jv+v6KiQUNl+B7hIHLk1Cir1Lk4DaQv1cfH+7qk1yJ
5yZ84Ju/xUs554ctIpYsBOQvB96PIfS8ze810MsvfXXXigNiQdRSQWYcbZ2E8m1N2vdd91IEWcwI
RMHJ9xWz+OJXc3hboEIcud6nQRBCbSXfxY2Cuz+wmaJBIW679qrcpL9TUNbRbnYKfkrPHX1hqygv
o4yYXj+eGL1U6MkF8Booe45oDBDF+IYF4V8dC8E6h6txatoDITS0I7JRASKpJq32Fz9pJqQweedW
/qJ/GnJwbRnacbt+QEaP2FjJMNnYIsOIYMWkk2kJU0hz6Fzwc/5TQ65YfVXghllX4be70w/+j7kK
Nwh5L3Mq9ExFrJCrB2uWmETKAGwG/tc9zm5AjWbTvkdTHm9ojqAGHe5wRnQ+fL/JsN9VZxTIyV57
IWbD+lSCTAJ7EArhigd1SKcmOJ+5MkBWPp6uwsT5DRwi4B8o0TZY+B4322V+lmPFjel3VyvCY7dh
nyUGGo/DCaM+pUBeXyB8eK1sndmOl4M7tS/V7DjEGJU+rlTRn7SUppNOgPWo4iYlh1d/D7vPJCIK
/n8jk/c8d+2AnF/ddDlRhOihLd5IhXlzrw4sdaFL7ClFOsVkHBOTRCNIpST5dYbkncDX6uAWYXO+
wL22YRH9k5hDxu1ud5j8m7ZNcIQqi1qh73dFxTAGp/hqqpmpBorrySsgHLVwkl2kbtVfa6SSK2n1
YEfV4tGEFnbPtSzFFSDVuE0SZ4CZjSBtxC8Rnu/LEkUa1cfnwD1pYAvcyjS0uKnMWxQPiGL3mXba
3AxvWZ2MiqlBma6/hYS1BvER5RFdIL16MZIrORUT4oVk+MeSRmF5LR69eVSfD/vKgrR+CTNvugou
ChfqTMcZDJQnPSNhE3BD3rC3TmXDe88i2GLYFFAvHTzflKY6OreqE295DkYJQW6rSFMi0SeG0+6z
y0yU0yJZsqEEsk7QRQxnMwJ0vcqF3Txyp/5DPiuEdb6k1PNDz0dGouOuAIBm+Ye/3ublPaSyn4Np
o9ZXI8q4CyZ/dfmvyeyLVP0MxoLnz/YOEu74fMhfeQvP7GUOCrgpuN7TGoQKtfzuzu8xuN8zBtdZ
4JogNeUhQv+fYXHS0ydyvcfloHCKgHKZ90JLkms/DzTej/KbwAyfOtsK7BEU9qLY4qbQK3Z7WLYe
7Pg+sDPqxy0CuqIPuMP2CJOd35tfzo86goetjJqCSBLaOnOi6E4XWDHQwgJKWlZuey4KMUZKLg5l
ItxFnVfuzypPmEaOTbyvE5de6q+cflH4crcp2DpMPQmrZns6OQ2NbLcfJXANTeJWFuKfKR+KDHeC
joaSkERsAPsNlXIsajtR4nLxoNgw3DBlNQ4Nr6Gr8sX91+kVmnaxNTrRD7qZ7Th1bvhVEnE4gTnb
hi8B7ScPWn1PdXe1E3SuBsqIoxhlMGa2wJBy+FFBHu+c+TqKJDt+vteXiMvrM5NQ/FcT7YTuu50+
E6FLy+rqEvt5ub3J//p3+RppZEfeeYxIuQH4tab/o/PC9ayTtx6mNzG+e0sj6jmvsF+Cn9dEcaV5
FhpIxmT4FYdk6O4+6mZd5D2wY+jLmE+WiKkOOXMAn6RHyojU3vA5bICZt9dM3d1le+JhWoDlJTRL
YhEJsyfDyUjBtTE50nsum0GGy3YU6nEXUkperBCnP7iVTqA8Y01utP93ICS2KiJwRzjBnLn+Ldk+
PLCUsjWSodDbP6e0tdo6bveZhsmdrdIbHYRkTKSoVPvzSQXif3W8a6+Sr+VmXBiGFhEt44ZDvbRA
zXeKC1n2+ZlolM8Bd2vVfVAwiqH8cKGPCkcdzowFmigyQSZVaPVPyV0WCxlbFsqtE9WghEkmpUBK
IdCroTm97NfzES8OsHAEIlg6GY2+37a/wGcmrZgQo17RYdkbjXgvSPozCsLrPUMAccXVu0Dk1RqP
Wv+WlyAe7uy5HcNY/BdC6BJ0AGZolA3twsJMp62/vp83kT2YQmEfAP3N137IwNrYViaMt7h+/7sd
LJXnPkX68Wi2HLe/1PCGCmDex1Zlni9T4D6Cd60c17cT3SKhn+8zKzSENN2xRD1vHyJqmAqzpxh4
Dga8FkXOhYQN/6LTE/SmlzMmhN6Wnnjpz/zqoxT0liARwBPWN6jBKX63qNk9uxfUoqBehg4hsDEX
//vb2h6UQtufirDE873dyMFeevD4o6eil1A5XXrWlQ5hBbRZkPiAK2ld3R2kknw7xGP7JAY7m78o
hVq4avVU5LiYApGWAKjuAX3BtkT1g8hQ9/o8L1RIj6vfV3+A1btCcQSnM2QEYzy/TWlBtyNJSUW7
LIRSfS7SZy/dyAzCFNX1cqPzbuM7kZpExCzFpBgnBGGuwtTQypgWjzuIK+hp2URhjQ6TQI2jWOuW
swf3z4GbMRnzYI8zjaTn5ThhrYPSXCKJyBOely7OaTwgOPxrbimEJZjwSjGN+8UexzDKBEgQGmC1
l5zzRce0SFkEDVFSawNImr2ePj0lCCNWsribQnY0+MGwfHJDafZbRUUi2gGVi/FO52gc1ZqDPhsU
EO0kzxU4BUduF/w+pmT4iTFxN/MjNV+K0weONqoJMuq3Ebb9bgCZJRT/dG/rc+AdVs2T8zKod8dD
PLdiqVlq6waG1FIjWAQgLFVsrWS8cWCJ/nPK5svAvyFKKZfmwgq9NFlFvvl84aXgFJTOWLdU3Cyc
wuSvyH0SImcX1bS3YsZ3umq/Xy6lJOExkibZp4spoPcNl9XPU1tOFggO+K/4UvAs6MWsDIO3GKe2
Cd5CuLlJqT0mlUIqRGRWt7cupQugB3kPJTTrfYBnaHZjCuWCDqVAgDJ2yzk20SjypLz3DI67pqXy
Ne8rbeYS5e1HgntAABb8jsFJW9wQQORT0jmXhGvDzmV88QMNCicDpRV3pP4s3Zo0M5aLfBapCDPS
reQKRgjr5w8pf9gxiztPnw6A4a6N6JgXJAjfaYzNaWNp9E2IveZ/xTwgYjMJhHVZKQ/QNLRWGfBt
sUa1NuFoy8ei3kiWP2pMlEN9DL79cQrjQULVIfq49okiEc995tvqreBC3vnsIAy0KBXTfA4/1sdR
meK57DHe0Q1cHfEguK2LnNGM3wWqvpPm60SRoK7RYvp5ty9xZS+Xj7MHdSeudmoqykZ2FaSQ9qxP
2R20wdzfAg68UAxB2HhBOK37pEpqq1FampfymYkvrWdjLClooubuSmpZCifj/Z6OVEPdYYm418gP
0TmOP5a5gTHgwrFVpUnLEgPgXzWmMgmQVDuY1TkH/ZD6cCdMJZP4inMFZe3vumk+LzyKQy9sV697
TEOlt6Y2tvVhCjg+2RMBFv6jS/4WnohE4vJv13DDtd+o8ZF5STyaV2ZHGitkyRUvzIzTIhjU6GGI
jPN4BnYoTiKCFvEjph384Thv91imhj+bHT6GaWlTB/ZdVX3JMM3qKuABA46tk9U2lkJpEIVCK3Hd
9vdI7GvH6+QfdA8gcTAwIjRa2U/zoUfERB9pXVdpoRYDlb5rZR7se4NBCIPzeqXR5NiWDBxAerk+
GXkTjjmHjk6K2F+mHYXMIgauGsbOQBgAhxBR1iqSwceX8R9FTmmISe99Svmq01pJklQ6kNYPAHC0
nzwMKPU1UNsGIK3TgnkxU4umzBCyhtUuhKJ08QlZrS6Oe8Hb1YOB8/I/v8XZofgK+FDOoVcg67mD
PmdYJz+uEDG/yi6NHiIQuVJkIy0zc9sbFAd7XRQ4L8z8AOwZPP53prnRMZIjZasjzQfQtiMu3qFI
+IwveIQ05Y90FRYesxmOAsMJNAVIoW9UYaaj+Cy/iA0JQc+E8bKNtt462osZ0dUtRpGLkS9Tf4rf
wSFCrfJbOkYzE9pADrTs37v7yVgEwbKCoFgPwuI3EMS7ZBKZDREZ6jfBDQJBN0cIQEqStpFQ6hCM
jYESD31aks3qYvCU9sjHt7hA1tE5F7ukeYOfVBGkYdHekcjJrx0bjlP1blojdFpmqad/L+SiypRA
AgdiUxu9J7dhPoCz+4X2vl+aVZimTAY+1Dc3FFAUMrdXWnLmmcwU6SQG1zTsSJT15lHauycrLgWf
7+PWw5zMTyl7Fg/5VoWWz5lOPB7AMV8SgP4snPWaz65nHQEvYC46rwsgWd0dDFapteBYdIttYvlm
YTDwTOQsiNDM2a3HPMl43Kgl2p2Kkm44qr0m/tpQOulTUWMFxuFl7Yf/M6X1813qIFcxg60+5q1M
sJXziO4NN0aJWy/NWnEyf1CVOC628x4DFJlbu0ULYC2fgcsmicoUOnNBtQ6LIX4BQO/SkGUAaWo1
94H3gGPLxiu827BuMPaObpUt8kl5MloWReT6fNj/04TN3WkornB2kcC3PV/Wk2sT5Ee6GIJYEfd8
07KJ6D8Ynv9qxE9EXK/wyuky2M2GD7n7Wc4cl7b09NF8RLEy82dMbZJ9gF9A9Q3EfqFsalOza06u
MvYv5xvxtTCQ9pgoyLf1QEcjS4l+/0lvvivLGJn4lIHn4I6qnNkNeFijVfKddCFdsc3TQr+AUdb8
AfKo5sCKBCnxjqcsmhtNjt4DMXU52C8EOSaqxQ2eDGeCYCM8EqGNLlqgcg/qed6ROpNtm+oILdnW
GAVFunF7KRLI0nBOeQYA1Fple8lfysWxhyNgXDwEic1dgBzUsxmDrmpWIWx4ZxYheTbm2xn3ZaaM
5eHh03ntQn5EoMTt3pz5qqTFKuAVRO79QvLPDPSav1BByT12YeXGGeMWXaXj09fnU9Zbwc0WckWg
13a6DPkGybdEm7N72+YYB5U9vUEggvTXJhNxLxcKdcbDHqW5hVoJzADUX3F0DiRJGnObqGn42o25
Tt/n1NLsa5u6PgVBilVmAgg9sqhwyvGcSGq7I3fYo0ceHTlG94kW2GKGk6hYT5kpiS6YNgpcBDzr
6zcjWSVdSYHXwMB60EdEWHYPUZgKlanrDWh3Lgsa49hi9KeCKwA6eXDm0AE7PvMB8feuWW75SKQk
ZLAL/mTmthL1b7AwnqLpZ0VJLmZ0XqxYZPzAqr2X2BuobxXnS1Ig10QI/6rtQG/HxG1Ss3xZ5QYh
I5Dj9/AJ4/rT8t9IrFynlRYxxZGJHyjOOAe/oXu6tHNHAh5URwbT+Zvp4bKcd425oEuFFvoux5Vf
oHbgnRxdUBgMm2wayXBZM5lht6uZb+MXbeTgTG0XCrqE2fJu23WWt1EEKWN8/2cOlkmBHV15vjC9
p8HE01JqA612gRxiM1PLREumpUpVjjMoovO1qP2T0thWLeiNdnxk+kweNQzYaFyeAKp5nTC1aXr8
tfnzI3Tkya1cZ5zoeEoJU1WPfUJwZCJ8VxyH19dOINmzvBADe01TZeGMTbSbRj3TbWWVcUXGlGKD
kNwT16Kwvt4rqXbQAnc4nGT57P7tfFlaQRWTihy1THzo1OUjGNuUPuJEIglfmvJXOZeP77/AbBNH
Ys9l9YBlDyMT04bgK7IvzBvkPA1FYnFjiAo5o/+QPV7NNMedZHD/1fRw/6jZbdnNo5hzZM2YwqRC
IJVs9tDEW8Yaw6pt+CVkBGk6zuEZ32TBDJ8qmNnavypAcez/GzzeyGOD3PLJSrIvoYLzxDkLtWwB
uVYwuNDnAoTuP4ZuBDBMJGrXlU3/R3iVfX+1Mgvd11o+MUtf0cBxycoLjE942jcXK5MG/uAMuZPE
PyTzINtCYaJ72ryk4NEjRWdmiodqVNP39YyhEe9ItvcWaCbmAYYDLZKS1ovEFT1rf+av7rMbMaAr
Q8TOkGBuiAbu37Iww+wB0O1n7Pu3ysAy4lrjbHcQ1PHxIW75L5mDOlsPHtUDEaLgfnsp36Ly9XlE
XEM5KdDxI7HAdVlU0PaBSs6oYgUX2YYYu2U/zV6erAhLXtPnzlU01bd8oOg3VoYtiGPSZCBF1bnH
2MHpMfFpkWrDV/4AFSQ/FiTiO6q1aBLel+oleephAjoEAI7reBGDOnwKgT9L02haBrrgh1xKyGGi
T3xHoCAzN9Y/cdfE7wAFwvi+mhmYl6+9Zdaqgl3G1i82F0Qve32mkNO7vT2cF7xh3SPUu6tYBfl/
2/12PatlUHEKckeLX+3y0/L2/NnjKfqePdAfwFC3RNSzglHF9AJDvO7SuPnEYV4JXKv8IsX3+MNn
lo8pmFqwBoZPSnPxhvVYMOvDUb5L2o7ZKbG38t9UTUPp7XCdJJd+br8akWrBVdpwvWEAp3FXOzHF
XzZHSls9BES1Elt9uL0U0ezozYevTMbh2f8OZCUvW6IYHnLU4dX6YwDulHFalZhYiRsbWoxqtYyD
mhK0ZNlU7PitMphkcTmWOyvpwaEQ1pjhypoCifbyycZ7EKqvCsL/eWvCp21JIlPWziEiH+4sXwIN
NOyIKrHI7+oRhj0xZ7/Xlh/DKHPpc6zqCXPQ/G7/DblR0N4tqSxW/EQeEpXxP5BetWXfd+WGT2Ib
YS9p/727ll3R8yGu0aYlG52LGFqk+e6WSI/HkZjAuhXtrg1aNrx3RIWgfMPP1PGQkAKePvPCLg0i
/kSWzuNO1u74D/vls+UlJthVn9fqsrbOxiQAW9XLE2LSM0wij1SUI8Q1lhgpmvMyfZOkJQ4+ErWm
KeokBDHOIL3UaNmzPU6kg7RJUI/3lsX0mMejaXj8pi4sEV+A90JtSzs1arE9j+ttL78jzN+FkNIP
lu0UMhtPGQ/zobQSpKSl01ANYZPhUcBS/lCQzDj1Y3Mbkl20no79C9kLMqyIDtbRYJB6lQTTirKv
ibOAan8rFQ05NJ5KMP4v2ogC70TBLamp1UMK/9R5VnE6ky4yEfgAuloL6PuUcqHeyPIQfCQiv8xS
8h5zTTBKdonXDfTYoFnP6AC1F3haC/VN0NEFy7rtvywzKfJP4qvfI3kG/zW3cDmy5YSc0kv3jNbD
Z9n69hflxQLvvoG8+l/p8ZtQiL7aWZb0qPFBfBjAdc0Co0rsar9KUy4zzXfuwaJm8BzzGL5cd6z8
HIaJ0Feg+XJca6zoS5+zSnJh8/647H26eHYMnt+/v7/XBJpNssFtb9j6HO6KsjtCTRyQwSvhNf0H
yO9bjGRhaXTuhRUhMHIL9XTZlJUwGaXymgu5IQOkDzNd2GzyVKbBkcpzXndtEEObQywm3nYrmG8T
b6mAHSG6YSKRNckEGIWpWtRGQ84RK1zjy44qxcEyTNFBqLdmG+/apjLXN7lc06nLl8TR+kdBtYAe
ztSlM6uZldMtWkWv356OMfg12asGyIAeShVRwSHqBmZtbbdkCroVCnUGoPPF/kWemZBHR2K67vJU
i/VasCgqFY3dMC5Dzz9LOz/JAmvp7Cx5G/PFnECEpu8OMVhj01h/h5VhwLU0Jv0LjGjR48VljM2x
2Zy2SQfHm6Xw1oqBfpD1i0c/zncA1FbzXGnHl4hFnC6HGWyRPT08Ol26788H86qvNICg+t/vLIrv
7N8+jB2Nn9Qat7vOxOAUz4b0QW//ifBrkn6z+A3PbDNmSDviQ/8395C0kF/y2cFfyaxovTZuFWyh
A9zPsiZXBHzp6n8fwgRKXiHEWCGbyWY52jZaqThjM2KIoG523kCoTm/zr+ULKJAEbwAu80WMGOqs
FCf823smledsLXJNMxDVx/L0CWox0ea8AN/kcKYNR4LVFnJiwe1Gk0A8xr6YIMMY/Wvyi90tRy0C
hRwpUlP+7kDgDTfKmY4Aik0CZWkiTiIAG+rGA8yJF3GL+CM9HiJP+RoONI88DIej/HfH3iKIkNJO
xRPKw4JpzOW2FgIAmsAVOlwsV8RcwPGEAA8wHYJJ08bPv+JzkLIgWIGfSy0KwapF3Cd9wVN1a02g
K9aBi5KiIhzl3+rBcxwvRhjSWxvTSMGBhvDNvqOVhD94bOS+21kbZ/2+9swVLK9IeAhCUMvt4SoQ
R/+TewpY4tw4wJFn26FlD/ArlTwJvhoLCvsAnk7SnTliplfaU1xon8wDHRObZ97mIcGZ1Am1h67L
yB2GDFgRfHmbYI9k8uoWDog1UQ9Y93OMcTGK5f151rZhJx8nBU3wAyMHmtrdSD4d1/jNK7Gp3PCh
R6bbFDEH222JNX5j/yKWXkmOAYAS1LJi3dJ3OJnZYgqfY4kuu2gSH30YvDieLCqulD/XFdwNgqKt
dvOB9bPM57nUMDRPZIIPZah8sjNieKk9GKrrU6CV5tnUAdRtxfoxUPhBCAYVckhVSakFq6JAQeur
9mfGAJJjcncPIH3261eV8ZKheERkDJsBFN1KJOdm+u6vf1vX5E/bwvE9q4QAhaARxOsYQ/HGGXHr
4ktGlwFmkoBrFCRvA7aMtqFWY7axPPa4C6Mhbh+qd7kC96B8rJpXPBNOSu6+0oeeysGo6ksvMZP1
cYcDYRDjcqhT417q1vb/eCZBWptiioeXlRHTxbDLAzx1Behcie7cO3+IvqotqOxhZ3qip6hpDSTk
9HLrWTp0SpwTUZWe2duWvx/MpL0RtGhUqQ0rBP1uaiF3CLmgPbhqqeZ1ht1Oes7sjXUsrHL/Tcin
VZbjdOeAVV7wjp1HhP18FnGfymasdLb0QCbiLOeZQjcE94hxTYNVTwg6fyMFW5UYnC3vY3y1/X32
y5nRPbPUQrdppUunMs1k3CzNS4oUkWXLQnxX+qQ2zEeuV1hyvRabHju1N7qgnpihw+Fs2VAt7Hcn
luYOnbNqT4TQjoeCGL7T06NeqlCizZLCrDoRGBjMLh2z8W8MmuTIMJ9nocdCEbj6CVPlrvOR9rTE
Pexcg+EESeIxNvadiyeejcAz7QZsN0v12G8XM4/OQeIsPWjzBoj89nN4f5m9ojWatqDqvihl6zJM
EfnXqzr0INjON5xv3UUjZarJ1pxlVrViMCUCQWGFNt7AYvgGuIlN/r3Ho61/EgYBYwj8ucgKEhqW
+5kSzm432W655VqA1W0aK9mSrljtLHCojjRSIrFi0YI+4lgQREav6qcEC4xgRzk86Q0sLgRnPFkH
N3r4N4viFyX12AWGo3nuRIXpRf9iQURCqTe6An+kIbWB0c8r5LS4kDlV+3ZfR4RxPVn+Mi6U3Pnq
Z1mRUBPQW/cWO7OaGMK/uk/Zff3mspyLxl27HsNgDeCgsy1ZyYdk2jiVVT5y3g3Lrlgqswx8JJZH
ZvpCYEJSRAY+YYZWJIXtTBrMAlyC99By/gparZcL/iFXaRyLIWI5e101o/jB5jeIKTB59V+BCXDu
G2yXGBpBRuxMZzoJYi4PJ6UxhK8HYa6IpGP00nHhBatiCYp/JSndPnmvbeSF6GIQ+yIyf4lKgbeD
w/FoGL7zWcR3lrXjGr1xftznSddf6GA1MLazL3NOmaI72uWv4WaJKp+qdlNBf5SFH0bJXMKowqV8
j9vMIYWd8nHa3rA0cnJ/ck5/1rLnRXmHjM6UAvj3VApVVj9K6xNYh0LkkQ+8id42SYALvGst0Z9V
vm7msGw+E91vGcn4KLzl7l1GJLahNAwn2mjyKs28NB915MVX7NPqJOtjoHC7Rwowq+ikh5evkAkm
tg1iDTo7DH0bua5GqDMkbcWQAB5CN9fZa3ZABUaCyEmuLlC0APQGmDDLXlKuB/sO0/rHrCVqkXpr
tD2u6kg7P6oiOJ7bWLzMbahAanLLGNQ6LfWQTsIJOaN2RWLfUWYIAODurjbbsAEVVMp8Zsah3zNg
8hSkvq88FcBl5mJCcFPpnlAXywzMyQPyvbzqguLjOddsLaaU7S5LUfx37oDY5HoTGopotIhQCC8t
JrvFdiUKikUgtt+dlulYIVac5NcFzlkiMLBw1boo/5Otux2iHp+vai6xgd1ZmHCSYCxTC5vv97yi
JvOFzBhLWrY/oOE7X4nZzRyFvq84i0tr8FeuETn3JFhcAQUNZvCZ8VxeDSf7NFGlEng7fjlHMzG7
MIDtnZrAAOY4HLydx6l8j2ezOD8lz9fyGNBcfSl+EcHfS0JTxOGAgWQQi2EJqX0a1Mx56yKhbELv
N8MWcboDolQd3POn/ULov3YdsKJ8dlYMgTSa6ySv9PX9ZqV7lyNtHyyNdducgaHUucO3G+dKP5Nc
2veMK+teoECKv4Ma+HCiDdP3uXdMC7Af3QbLAs7eYVdgd2iAZ9L7EExFWULn9ETJrkAa17fG4qi5
8Na6sD5t9pApBt8Njy8W6B7L/qEK6dUno5QsZ61U5rFMIZTAO3ibliDWnzYPaF0gXyYIno7RYnzg
sgHYonlWFSFZHi8x2N0VJ5+OtI6GEJyPc2ScxzUJUTRaiKV0jj6tBVQZtWvibBN9AkrfQE3QrPbg
xsIQ6A/cSdg4igBVOi10u2tIsT1HFXrUHY0ollXm2koXqakPU0vaXZRPzzGYlGQwRKn1xSEe5Xuu
SJ6vSSlWlaHKHoMxNy5gBZ7mxoxMfOwEScAKSCQ0JcBUj7j5RDb/p5UUnvrw7HHW+gB7DNhf/LcJ
eszVUtZkUe8zrttspR44lO48Et+tvYvZrn4xbQUNonsJarkk4ZIdaggaOL+c+vJNgUQ098/UoTSM
FFOGistNtG3p0Yz/qhs+o9e/C+FbBRYZo+ncVB4AhERN/NrQgzoCE/AXi16Qwo1bVDbicx3GCe/i
xr/J3/gnHueJs7k2h4GJpCpx3h1kyY6Pttsmq0vGnYL1f/0+O6eKVi4bVzAtpfzF8PnvGgF7HxGO
3eRw5/2M5jEG8YRzG8AETIiS7JgcWnGREV8rRhyIpFEDI5cytfYfULW6R1wP0QBgJjkF8I9wwONU
H0MiVbKypekQfy0cofXWKxwHdKoPmqohM/XcB3q7FMI7x5KW+LwIVGCmgdL059XpEJ7q4iYdL1o4
60jQol9BULNhe/rIT5kiMkjR0o6z52zNGqN75RQ4N4FyFhqPt9r8RdTADLemMqzWCTO6/WbArvMj
UlNmwq3sOpcEMg+gtLfIJCfGn7/IHKHBvvp3P9mBoRG3FVid0ZnLi5A0ns1+yQ+i9H8NmmQiDOF4
GV+qqcYx4UOznLbWn5sXIerU4fiA40u5fnviGpqGLczBY0JH0dCWetKMNOn4BopoJO5PB10OZsYM
eOjsWo3XJ6OhvwkqKw/8qX8faZeMJhmzJ2O1ZW4XmJghdRx4TZcv4Pcg+8gNAxrUQDDYiwVldkmJ
V0tJQHgyKm1UzEPiNI+DKNltJDbZdq6KoyrvapEMZtlqzEi3qW8SEsRCxNh8qAj0P5aov+1EdIdH
cVKw1ncK+rNUxDoREgpV0qZg3IEzuJrrDE4t5f0e7sR5ct2DHXq9LoHc8cp1juEf92V9KaZbih4u
GcIfUuIEwu4RH0IdZly5nH8KYp0Aw5crZqIpOINWQu+N9m31XSLbKt+L1QqO0R/KAY1V1oI1P2/g
5HSfoZLWJoPBWya4Zv7Z4KyAMUXKWEXips/wA2fXMKKdQy+loIIHHrjt9j8HIrJ4rl22m1S8999R
WwT1s/MgUKpPEMQG73tTe/2cU6qlfMZgVIiwALHQ5JZOoccJX37uybd11kTYauV3A7qvS1BKSYmE
y3qr4CT/dpOaj/O7iZbR9vJD/dkN+P+VRdE+/rl3j8idoU34jKhwA+UL/zxNSq1aogNgigo5MroD
LAEjgIcnSgG4BmPsaM6UzqWi0zU+DMpFmsHdYzBVQUmml2kMhJj3uukJ/+C2zmvxJvk6wf100+XR
LSqfTDSFiCFAzv9ygrZ7Xb2yUeD4B+SdbFil2XyBVd3+p7xdr6Ygm3M5PwkOEy9cW7Akn9yXg+4w
H05jcAsHboTqWlmygF+urKz+rXK7/Z8KhX2AHzZ4+u/70A4rUq5n+yVgYTbXY4v7VoFdGzCjHvqD
GrfaVW9JVReda1GDCEbNGd83VPRzC5+EPa21bMYKuYCyyjevqJeoUP74SKFeClJSdhchYHQrw/1I
TpAyptO9MG75qZrZGzpWsAVq7/Hi0AiKembP4ZzXmeuCeXi3ySm8a2nMlzA4JK8UJ50BXLBceV9u
p0PpIbqjZR2h36ssX2l5dHJUeNS+xNzDbUJKGIALf7X9FNZOKIwJ7j7Y96MkI8pkJroWXQNluSxs
XWWncmcwpCL3iFwB42hgF11QcEpvDa6hBU4Nw1hojYmq8Vf3Tuk862uCy5yin53aPMNcPbMz1j7E
MVAPt7KSb9UbgptlzBY/yAqT2xUn6avHWm27935B1G2EhUAlIJXRmeieZp1zEJKUH2t3f2kMpeHx
d+MWDvvUDY3yExkO6wccSBeDYzJklkKX60m0dpYE41Z9LsqYAmsmXFJxyHUuPopPT1MN3lEyvz8Z
UHf7L+t0rMdm+Us8BbXAG3ClDQRW7fdoTd/bARQwf2yeGjRqtlTk28Yk11qBOKyILJayivjhDJUm
iLy8UlRcIsXD/WZWhBlkp+C+MULbs0XODccZ3VhXtDPhKQUMPq1oEFfN08WdKT6eEz3cI3lPu37S
viGV00AEee0I050yYng4zK3UDyd65sxB/8NgfkRnUxXCAacef51Cq9OkxMAv55U+JnvdMVuniHWd
aONSH1mAJte+pplp1GHZjDVHuBJol3FoEaq3aMcAhM80JVevmH0jGgRz0cq0IoTR1L7g6UGDH3sg
V4cksZjUUQCkbd/zX5C2xQ8dElbhlpJGWqsg63RXBhBIu6nNnPBF5k0D89nMt1RDILhFG241v+F8
SLgAybcq22qCTt1MTeK8UJ/H++jWttcOJm5/AP6QMOYTAKt0lhHQEmg84djgHuWt24E68jmuvLQ6
gZHVDMWjUbg599Uz3Z5fVzydUhd6F5soCXcNmj8smOfoQZx2lITh3JAv9jrJ8c62Myk+DJKy+YLM
kd5dihDeTvIgv6p7NBewZlC7dDx/r4YSSzb7WSqvl7PqJVt6M1hVEyy2kOF2Ml0jMcth2jNvdDtv
t8sp5qfApWw9ALupBpnmY8PpD899wLhdRcZAuELtGkCzz06vNKrhs5UmaAuM6Fqe1ntJXwt6mueQ
IbmN3yrzuS4zgYztzEipIg09c0VfAbaNtf9RhijIztB0XoML4UkeniChJvWciIOGLim0Y0bGYurc
3OX5rf43Tkhh8xyl/9aNCF/7MdSVa5rD0G34Rvkc0B8fW2y6g+rvZ+CFFTIQW/JIA7WVNqlmp6+C
mk5ZVeAQ+6WAukuU1gGbod7vZOFTyHGx2J7XuVj9sr5wwAD4LwvWwsEFw2U7sNCrLNlL6p4yJag5
w+o1MIsgadHaDh7hnk4VQVY+kslMKya8EOKtEcyKrQ1Tr9jOG0uWDposewCMgpG5vX6ZIrOKPS/K
syjhvRMKkteHznowesBQDOblsTrMHG2QolQAlF/W23gjB56is7/7WquBfhH2Dj0GN0/TR59kbP+a
CL8t8RcFFu4wnD/FsKXzXAqBUP7wPws15xLsloJ89lD+q/7uKObTzf+shTXsM354teHeMjFMDXSl
jxPeaoypygPo4j0yrLSYsafrO1gOxBndcegj/4vuAIqsrTBv7WKF6xlpRhusxAV+o76z/XCvmlw7
iU5YuJaqC8Pl/JGCEEOLLqhbNog6rnSdKbX1kby5yLmACahJmYnSn8QEGMc6gNrJMjXa1xEplVD1
tt3Oq+ALQ4XrQPXxcdpsyJwwsONFklMGoLUGycS61PzAjMviy8BjStAz3ZBUXCMMfuso7ZKxC8V0
GgwQu7Dte5r72wjsInEMEi/rMopFWe+fALabNApxwH0CT7BRGLh6s4anQtCKCgAz0wnd8SARz0+3
xWXyx1M8Z7ohjgoFmNuHuTOdAxHPtghUWkigRLG97X5MTiFWtau8TO29XBrru63mM8Q4sYVQ9dmj
8B3919/UIAh1spkAtiFr4oa7NL72Yw8j0rYZA140Cyf4jxs1iMO4s7VHUZyy+e5n/cz7kcDLS28j
Zm6kZwJjxc7HFVKaT5EC6MGFhXQUPfppo66o2LDBqtWk9mZQPOEvTatPyl8L1gJ3uiUhcnDsynFM
4X0NcxI7yDhoXsKcVWvGMwBBKlwCW21IE0wQH99GNt7jfFhSJFJ/DYg14DGD9gmWhHOZUEBpCnJu
gs8QqG/aQG3yed3GCCsT1x2PN2ntnpF2VVI0xp18YA+BYg4sh8nQfIeB6akp0/K/V1D9uMpPancQ
WxK/PKFpsmjs0drZ0Qdo7V5Yp+1dlVCKzAQObDVUInoe9RgA4HOmOhdWSSnG/ZVtZ79FCJulSW7N
t4hyJqulAjr0NBtFtnCcwXJPoha0PaDU+MZuP28QJJlP3SVMgxf6QBcEWgpLyROGZo/CQ5oltki2
41j3GoUXZTcrW7WtoZU0VSSgh4d6k4NIXFaeCR7SQN80ksN1SIi+mrON7GN2WK1M3Mj+h8Tdkd5H
MTjmhlMHSZ7MOXu8f7nmZPh9bD6SI+HURySg80F4VTKSGlAsoCyhw6rYnWoPa3k9XihkupoxtP8i
0nse0py9ANm/1LMC9EYUE8TjNfY7QKUTJsqntdALX+E8zptW9TNkG++b0fnsKp2TJVNty0C3vHJu
mKlgUZP8trAJQxDaHNcnVy0rla3AnrPUGQhdDPKuXqP+o26CektlI9rAQnXD+rBv/XquCZAWZZVX
dZiDrO5rVtVPunVkUAl86BJEa6QUg1BQQV60UYAjDqwmku00/pq+3xL5A7qrZFkhb04fWIxXRnkU
MOQEFySpNoejVSArqyau2YU2/sInRQL+RVJgzLtJgL3pJ69+nTrAlcI/Br2QC/sUhC6YVBQrAfyB
mml2UTXgx3bH7PauSdfR95xC0ghChI5n73Zi3NOMCZ48b281RNOSjm2B9pY0efiCrgmLy9b0kYex
R0Z7g0KC6NwfwDUectBnePC1LxTbZn/nF9+6X/4WAs8DF+P1jEwRDQeLN6hRfwjsyYNh/Jm1Md/+
ijikmDixcDAkag1oC5eeEAC7HYBmqC2Lz7KlShx64tlyMvsJQAzQUEhpHzDU5Xi7JFwz0nrT7ROj
z8wCdm25cI05/TSWPNslFH3baua6oyfJHkkGcBiUy845HsmnBJrAQK9VP4flnN+DsoMpk86SHImV
D3vGhdH2JZSqkdblMWg/LI27+17GjT3+F7xhCpiExNm1UfDGtaIV3jD0GGBxMop5ynMaQPP50BGG
XwV1uJd9JzSnjRL6Z9t6/bs2KScdT7hLGm+ZZXO6odtIxv0DzFyBzxOGkSQaMaVhW56hkcuwGieq
zlbmQ0S3c0CxBxtOV7fUi0e/RAYh8pe4DdCQRbxAE3r7759Xxx5tpmZckI3vqIsb0VySqKtFy6d0
Peu8o/cYlw32z+T2iuPhaAAq8vw95Px72zYnu77DOPqAjoXpFp8dBem9zJx8pNjdJXtwWH9sRn/o
4dWjvhInBSxwXdy3RTcmIwwfw+ALi1HuvBg3rY/QPsz0dD8uoJt+1fvRBfcEzPsk7h7I2cRe6Nlk
I7fzzBc6vH7APvz3io0VLSUs+51EsBOYJRa4wU2aLeVn3DudIOp40XE/nZ6NBzhHPhDBnUdEv0Ok
nsBySHnQof3OCJFJvkkwtcw4icP9MXkyWNqLeaxq0tSGwKBc4MJvOtsx2SppwO6/KFqwmi2xXimn
AasH+vpZgqERvthwlBV2i7ojHyTpVfHQsG+P4XsxY8QnbOqJugITapJRF7b/JeO2n0Uu7jrzGOrv
Qsa3Kn2OppuwswO2gF117mPqWqb0NBVgLpQOMgXBYeADSJu7kexymQDBSlaPM6aryDUqOfUbPgTL
lTy3pehIyj+QBJqF4zxJ9a+b3h7qnPwNRAUUvZJpz/hfrn1LeaDREw7PkT66VpshXXAhE8MKdsoY
omHvEMObX7+Oxwsxd6QBPv2tyRKBJ9bRV+CjpaY+7jLwpkKmoXa1PNecUHdetEupHbEUP8N7849R
NTRVdLppL4sYPRAIrKDYUE1j/jnmS8fFNPeDxvnDBzFoNVMNzvL3NubUubx0QdV2VwNGxzn+zAqJ
MMUSYuIBuy58Ty6/H8hDQm2xmBkd+JIxle9Zt1XJSsXCBQBmHuOgZKc9LGZK7Z2/kEj0FK6/tbv4
k+CjBx3qtsZEOa2zK0yhRRoiE5zzPSnyFzHrQm9F8ngLIOIqAgiqP1FPVLwykZyft2pcLitmQvqR
3be1hXYSg+iC1Q71CGWYnoVwBygnMoOxzU0IUg2BBWj4xeWX4Tu2r/ZtUIrh0IXrFj7LVXp7jQ5T
1/G2bVp/mWCy4Imr6Smn0tpcAibfelBVwroZ7uTGMaSrEmz8ovKwtS3VidrzUCrjgBD9uJ7TpFbQ
d5u+RcDuZKkM0bKa0lL7wq0TyoB8upv7ubo7TDOh3DQXTjuJKRfxUPQGkjqu0y4GREAkayDVz/Qn
B0Tcfb2o6KDay6CbG/zNdlxcdkyP0jq+YBE/kpTDNyNM0cJO5+q0zP3N2pw0ivNbhPUeH7Apocq2
x0J0Kj3NqUfkuhQlNcec811fkPrzhKBIIRYFTt77xL+BttiwuJoUOJkJWQQ4wuhmGU+nFeEo0thk
h1XtlG89r1+/d9IgFTA7lX+wJVVeRvQtjleC0M8TH1rhjzfWAu0hZK44KOnb7+16JB43xriDWjd5
1mjq+epEjXz4WA0lNDPeD3cbx2564KyvjaWI7fDGZRGxQ9LwN+X2YveQra21Vde9B+Z7XMQhHLGp
dX6afuM5hr7fd/t7X6NXcYoVgJVFFI40iBv+R6TK4W+JivoQz2C3tvYZ6u8psA5zzRSsOFZ4gmSN
kBEpHyViv6ov5EonOyQfKyPFIOOU/DHp4Wp2vpFla+4A7M31u0M5HSw6BhYWIlVq1yFbD0lJY4XI
0jCYhbgLkfap1VzKr1S+QQ3vBLfzoDEPPOlCQPuwZLTrQjpP6zraIdFlz1ua10i+GfiJT+62BjpI
/ypJ7OE9sx9QMcsug1Bw4B6ZhgQ/jCtGXP4hxqwocdAT9C7LsjH5+wFS8HfOQcGIafWK5hI7CKLx
wGLN/cLUQ0v5eLbPRPEtnGo3vu5iFOQK/IsafI0z9e5RKC23cwg1xYpFqJjToUKfUgO3nCNoAtkl
wTh/4TyfhFp8+HFqYSJJsayx6ytDySQH2n/d/12exk3G0PDximRMiNxP9wyGwAm6f96VK3mGBj77
xEgeifAUOV6Hwbzm53ytaK7MGPrSFPM6eHbPVpE1fznteJYCPNIZ/RXQptAhoF9UmwFRC9LiEFEu
TSiVWlCPjqxwZ/c1qv2FWAdYaqjt8/qf1kUMSyJlIeDeuhbE3xBej9DL32BWvBCrqixIunKGdQ5e
LQnxyD6seMg5CmDrwOIGg8ek0pV6bnSSnPkVJVwdhdIhA55yc3QDDCQrmlcb0lfxtq6Hfhi+YXuy
i8qjMBw1AOIA4WEJsTLICqUJ/OMZXOjQgHbao9u6HGGkVeE1JCcAoWZw1tOSXgU4nSgbBWv9f7IX
OVZmJREEwd+VYulxKPSyvoEA4X/5Wq3C2SMtAtJmbcJxr158l3mijw0IGk5+JZLMk0bI6ptErfUR
df2fStIeSd72zTeRyfCY1+j9Yq6OS/PeBTF+bwQxMNWznH6ughCI5+WUXBGCOiF17hfQkkIyP/jo
b9yhzHnHmsPY3Jiv6NXNbHNocUOOTwWELx9t1V58iCT+oNXAEu1iwnWSWLBy4wkoPrkMj5aBEHa6
tXev4OvUQWA+N1F45uEXEXynZEZv1/hME/gpr8Qf/K1WXOOGOzYTN19hXXAYjApzhna1AEcTF80C
Wiq5HACSTza8CZ+zzeUmgbf0wt2ai3UUB+zrwnkZqZoRHm8DJ6pqsceJ2XPdODTP/DyPL0OS+99l
ssS1ZHtwGZ5/zrKI619D+xTI6NrQZMITIbEuObueB8KcvyAKrMus/g7IOcZIMKSfN/4V4IkNM+dt
/K38m2BhMB13sKm/+eD2L0KZ+OxJQqCi74NcQnVamC/vV9hb75pUPCMguZMPGe1AcuhgsQH1uNh1
cxjBvL3AuaBMukk35qevAiC7SwxvNs/Bb5woBNq4PkS1TjprQW6XQ9CIaZ2v/jAGw+NquzDCjRLa
WhDqpL8Cf4saRDdf5DYT+cSjWZBHp0IgRSJv+1WEPONl6RAen+sTbaWCvfrUuhANbGKUF/Yq9amj
++m8giY1iMW9xnVNY9ip0HLi1cXnhMkQQSZQYipkQzAOxy0XdXAbTPmv2zlYBZGzYYXROML3bGUm
kJCU6nELDYKr2QPJEw6OfoEn84e9MwK5tEgXQ8qt9v/GGotbhfKeWD6+b8SUtEXh/5J3hr86JhoO
jZs5VeW7xMQ4AsI00VaBAf2KSiLcGmExVbgGQF1EEbJL6ssddvVZhXPXUoriw/dQNTbeZZTUBtfD
LPIrjETTxNff7aNz9nrF03JibaOVv1xVR/z0pTKYvz/8s9oUwQ+hEiQCoojSI9H2hFQNSm1SnALv
bH6MeWb+cAVyNyZHIZTfan4lSpuwieFNOVR8k6ESdFHGG5RPNlsHVdi/LjWjcHPuAPAlcIC/Ueq/
xgm4HlgVwq7YR+D5g+fcFky7NnTqZNYKqGhz8Ysc6evMSQR0FJIM2j+WElKnKlOUaBJ4Jm4jbieI
pOP7V0q4Go019Jtmtr2jCKNxKPHuGT0yt1efnchlqSN+asdjgY0ETIqTSjMww4F9B3DoEZSZPAUR
dDdD7R8YqnudPdI4/OqdpcEWJVx8UF0/LiIWYiZ6aT3U6ku5wJXZx/CQamnhgOR53RTjqfp8yCGK
mKxH+NDT4G6Fs1b245ZEQ4SB7tutN8TTe28B7wGwJDD/sRI8ddwWQlsAnDV3Qq9LnXtEQeGc0R0g
UCifG0VEgnaQ89dEh9ORog7MtaA6B1QGbyq9B9BfL1vsvdF4xSCpJ7z7kj+9LmN69+5j/KCMzSMZ
WniHgjbMgWqjizsNJU5uHPUWG8y6zEafn08QGzDL8ctowJbNyI8HBLfIdte741fYT16ELwr7Pifm
KDoLDuD9+fDLtyuUflwPjaooabh8x/emdMfNAILu5WxMFKxrTi9Lnv0VsTfZvLs937DWh8fb8vIa
xQ8HC5GmZRLJtBiSpj6Rl2wGakNIeCO9Mnyyc6fnGbLGfGbznpKcI255njm7FTsYOy/95K3texj/
nTgWo5jgcqzAP5EIpU1tIs888v1VYFSI0olkFhrTLlWk9x2T1WpY53o0eGe+gGOk6otmbQ0KaEAu
ZkKW7JcEwSOUHQgnsLsj4NoKbKHkGWr3XI/MH+vjSvpOK8MmFWS295MVc8PW/FUpg88ek6JYxFzo
KDWthRdba+5EWvzl17l0UA+qzLOZ0yrP3aY0H1T+antR902ih1e5F08OZJv5Kq8LUNjaV0Zi3F6u
ryamHfgYfiAwSxk80OsytZZHkYkLOs5ZsZM6txnZ3s3aHedzxCqPTxgIL8aD0dT+ZSakZ33XXxcn
Ha7uA5ksUssyhGomw2rFUdLCWa/fNsbQBIIb1lN7LbMipFaJ7d6sii8kPFpsNfNGYfAklV7nDn81
rr+W6+onYXhubcrdhoEl3O4CcztDXtfzK6XM2dgV1rcRvTMAmC/NmyFQ1929zdHoMTE+AqdNjEw0
wapFXe2zecBZegZhOHd6oHz7ROV2aQrePF4n+yNVBtKB32Yxi6Zd5/mcNPHwppr71XhletfdabUH
oBh4O0xo5ggSj/ah03clQ0Pru0aASiuQA4oe0hF919kJ7slj+BzZmWCUfH9lXCPjl2XuFTm9Msx8
6Z3LdCTXhs5gdjt9R59wEkrttvyIV1qjpxCCgoW7T9xR7nEgOkfXU1KdqvSGMtNNNErB5YygdRtt
+YFyZVSp68UzpqMHD7kPap7P/JcFNUPJLD4dYhk4amGguFgLob0Ga5lKRMul/Oc/Uv5ULQFvJCmz
m0pVZDBjLnDdflU9DZejA2EFO1o/wXt5BAwONoT2drhe/jMbbADZPDTze7jTp/WjQaOL7Y+EnUP5
f0RLFzkByDMKngoqnJO533lqrofFZ4YPauSX+VPCH3rDMvtibcTfB0WtmmdOqsm3Q46BY4qndaYJ
GwGEXdLMm7OjEZLIszZ3CfiFYHWh+4/vpswHb1cOlPLYpX8G+ceO+eJ0wL5UUXbVC/rEYB05ZDgC
XENOqaOoAJrqGO8etjvb+1dvFZrx9d/U+kKt9BiLgi34ocOOwWw/NOdMY7NBJa9SiUfs6Fv5HLFl
IVUQNZCzbLiSc49lXYcX5fZpJ0QRFwh3Yei7dfss8k4XRvIzI5fip31XsRJujG05hefmCJINj9AQ
klTJ2Nt6TZD7RMZYM9AOTOPGJFCJHrT5nHZLQxB8y0+VrFd288HqI5BZwaR4hSSstcdHyFFvf2v1
EIaCvH7PY9Jyb6LT8xwADUif9Ae3rtffBCaUtVMGek+LJ/OBej15/MebA1kQpAzEcYKyohTTuePt
2b+Gr9VfJiQDHslQOumNhSwy3QIWf3OQ3fNEkcZcsE/Gd31y9FycATQ3t2sxiX/4Jk1CfI7FXdSX
4NMebSyoeb9k2YMS7s7JioSZ8hOIDUDfwFjXQA2mKAG9k1JpiJQXrYCkJibhTE/21V9Vc2PMyd8P
my12xM0hIePJ5QO5hH0EdHA6lh5aYzpGRGfU556BUfspfB3POCixzfMQ+L24zlMAAMG6736btTRZ
e/5yK6Njjb+v1yQETnXH8oR8JRPmPyimnrnLMbVMHxZiR+swM2kD2Wf+evBoS43pcXzHkq6G6sAO
i8SdQlFyPP0GbfbuX4+VzSLhNEjDIi/2o4VfXUOnLRJs0XGqvRiVR0DcqpHnZ4tyuwm5498Z00CK
gNUov1O7MBbBFHuTlY0aaQ4Y4GaOR0Awzf0Em1VL+20okSCDN+6oK9ujrov2IXfLaecYvlf+C+QJ
CTkRhpU/zy1vbHKP+5Qb6q/7YUdE000PXmEi8tOwKtvx7B/at45ltO6xzyI7lAaJPIYorsSzT39C
Ry5ZzTOXP6cKGNeMl4Qe+YsJz1Rgcyfb6Z2/lrkZTFyxt6nA4pBHwJspN2dj+8ZZPZqGmqQsL/E3
064n8Y3LBZvbc/X9RJUg02bcAKaVB5tkyWhysoMW8+87B+Du3gSu4RtT/Th8TtI8krzq7Locvcab
CjgX+SKydTSINjbf2WD1pphXNzdY10M4rqCfX08fkWvp0XVwxP71BuLv0ZDNJM6dv0dR7e7Fa7HQ
ODQnDME6CYOaNmuvT2UKAgh9wEOinnZlb6CJZIh/WWtd7/EKf0QoAMn6TJrmC+QsUMBUj0lmpgZQ
acYT03knOLgHRc9sY1Nd3zjF17a5WmGx7a7YHi+Nx3N/vwxjBrSR7HGYUOFUEOEl9svldMpMGSgo
pKPQwPssc6p//P1fVimKqPXhWuCyQLDGmA2u5ZQ0+H77fR3TAweQq3fvmw0wEYXsHBIrdsABapql
QuiBeXpw2gOqsEi5rzJDyhT0MWIRWSrhuNiiOWQPd17VdVc+9VGnVfSvtsnd9rqcUATusu1tNkwe
gCWHry5yoAm863hb6iWyJ/SUI10JMU72bcaVB8y8xF1XmJrqmsLVcSocDh6LFAiQ6Lf6LaxQTT7R
5ATlA0U8x7Hw84tfEbteL3GQb8xaKlyp8D6JXeCw1T+Ym7hiwtVPO0ZE6gXXlgEgfM2uQZkMW4Kv
Q+CJFdq1bxR3KgiusDF48AIVOQb/Bqit3MW9GBs8SSDBj1swc8NkvgbyIHE48JFo4MeCTthYM7vm
T8IxWLn/IW80Z1Mf3crPrrR9TJuQBOMgjimtc8lLrdEC/1XFturR9+hniJb2AenvH8LVp3LixkCC
1hINPz0Bo1sD/7JwFZrEMQdfiRuD2QQOZfC8bfgNAXMObxr6a7PorSDcZq/xPNTTHQdx5yQha6Td
CS1occZIG1wCk156csY4P+TW01X8EyEWSf4pqZlOqKgsr0RLfG4674NwzXn4mJdPsmXerdHEYG+w
P3BP9zOfh8oYfz8+kELi11JLcaRy5YTmLSjeejm1WdCDsvljAmCUytorbkGm48+/MOZemKNuwq20
qajg8J15bfFUpxr51LFQ9GkJhrfIwwZ3Xume6cCURcCtOTjmD8k12+N9Tq9W4fvf1+UuG98/TflU
ET75Z6MySHflOcut6UZeJca+sr4GoK3YPhNFVtfvC6D6NVBi9wh0cvb1nf7UTneGb0Ygj0EyegAE
kop0Lwytxmqdo3/pJggOm8YatdJxnk7DqVwWpoNN/czmpXuovY15gqrKxoKUlM97DA6Y6c16Yk0P
cV2d87RCU+hOVq5XilzSc41qd8BfScRVgFNdVWduyIuxrzLeJ6roKmzTL8gVHI2c24/HJqpv09CM
hHksOQxRyJsUFCxLdq0FiLMxDoeTGEqgZVtPpGnzZsx6jWceqLlr/moVpCugjgidFWOaPxcKNtkQ
xvpLQLyGmztEXKnyq+BjcI5zHDrbklX0EOZ8v+Nx9d0UvM528tOtWP9A1wajiZbRUSw2IRm3AhAQ
gOdbpwerKf8g4eagRGfrye51Gw96o/3d3VeSZ7sD/6tnWMov8pmrLMWahs4/pu6Wmu6JKwhM309U
Mx4fQTUczUioDh7bPGCszezy9RTI/0M+fWsj773uklA1LIRDSzUesNYw4JWVLk7myHudc31KpWFL
3jQsMUfYKzo2tugilF9KQmEepZj8bW5JhGRzIn7iQ+WmrdV0/YTCkzDWO+8xPW5jRfLuaxrTae2O
HyT/C474Afwxji+XaTJVv6yH3t5ClwAj6uun102qWOsNAjEdDZl8ZnGBxTPqs0/shBducjlIIW+3
rFKHlIpohO+yvcmgQz+G1Gny0fhgTGiscQhGct66MG2za6rrHXLBjvZprd9p7PLoSTDJOXHS24uX
TNpTQI4ehH7MGEMuwzsQ+IsQ2WiKl+G3d7hoUDYveGzgREjqsXNxYBxFNd6NtZygdAnsX1WmGxPo
x4noBeFCwM4u+6vhxLOIN0yvHMZmFEeaSF3icloLgp9ZjY+FCpElLuInlQhoTOUjsY9IkAL8wip0
azcw/rC75guRevntAuliaTBBSypnc7flupJc35sK2Af8P+5Sj5oe0vAMf3WuZTVgMiEkE/NjreKC
6a5VC1+OWSbyO4bRVActsrRs/dZeoDi3GMiRkw1gLB4MFd145aTgDEzy2KNwB6FdrnnqpRiA+EDu
qEtw/XHj6qYgMLcnbinunmwk9eEmgiMN2O36D37gOKfY5on8aIqtOKMJbjcpYn+KLY4uN6VfwsQu
lCo+1GaaenRZZ2vTOhXrPU+1BaE92lFD5e96Oc1KMQfSpx7dYMjJ7YfQaJJq/bogtM1GVcvP2LXT
DBOsPWfjjBxM5/tcClqQmZ2XQMAXGr3sbDLQhE6mMtPHqS4qyEzfjXer8Fr6oXyu3eSDzfOKUt2D
NA2IQ2kaszI4wl4Zi6fd4vPe9dZjak2TncHsRnUzX/r6Jq11w2fg1DdpaXtoNlgRPeziqoVXqWU6
zaYJXNvcIPaSEcOEiPvyN/8ocSsaBDrn1qP8gYOIJyTd/27NO1JZW/EqTLUpD6vKEfFIAgZzcFUd
0CMjhQ0O3sFQ/qSbm+jJJRrIHzCBbGmpjAPQFAPm55oBpcRIm74FrXONTsgf5psf/gyWhcJWPPO9
0UIn+3ZxVkhAtL2srdKep5O+M2Rgv1H8V+0qIS8VcrXMPfoSLQE6hVDR1ziZfP6SfWrKmycuwyyq
FDviWgID2jUknFndQkQDJxKAuJYrgx0Ie0v9f9Xbo9yg4h+PPmVMwRQKAH9Eg0+SEayZBfXghmt7
7g88SAKRIlN2Yzc5bXYe26e7TVJtNMXxOLPmwR3cyB9NAcehLPUJXmQzWtrjyVkMNVtD2ynALS6Z
YakE06D9OQ7WzPQLFzIWiXn6TWHICLBpKxlboMcLQYbknh8rPtzEoG0ZeY1GF4bIBpt4UQRerD65
lXZ+rHcWe9U0CppqJzL9m5En7SEisLnRdkUaXGCD9DQgDBxks/5c5SvoX8AxGkG8jYilst9Xif54
GPgUDKTf0yiFqDfLt1TMlEIKe8iVldGM2OIVzP32eTYs2Tc7aRICWxXf1B1Lr0RLXuMkLZVngxHN
2BmLCLZSjjaNbMs65v99xqHrxK8aPDG0ibz2SP0GOe+JIoIpEmBPxnWt5NqLd4q0XEQjyGdTEvpq
Q6+Zz4owpA/yHuv3sT6qTI5EhYp4cY19fIu3M0nhxMk4bACRqKLMkwmtQKCfMPX1e6BE37AWqlGt
3oifbUpBxpXyCyTeDGyshaGXvSLekZlLImjKi6dSrrL/XuFKyYGZ4QsG24o3Y55Gn6SgFil6ZfbW
04Wvo0QBkIegJDm/o93SU4H0hfviJuE8Y+S7exPJCwdpGMFoeYFA089DnOUAf6axLcsTzbL683FG
wQKHWCu36BRDLmO06W1fpONFuY+oAxZQax+RkiAsBLHJjPaylmuTsKqHs18Em6iIs/hqUrfPOGmI
C13VOXrHzEOOLIrHCKd4PfuogRrUw5ziIB/2s3uSsWhgzJ4nnISyoR8Ca3qUBkSTK3De1t+3+R/a
WEwHVXPpmzHkg7QVAul9xsTDY/Usa+0lu1FDRsQ/tn4B3FpEwbKIbJGp9M1KQsbX/0B4Ix+hokKs
VlwO9qjqAeZ/oXQGNjlRPYN9VeZWMUlnnLTz8XptH1tAx/gRjy74QmETGHWe/gm6ownEPNBeMcUG
p2Xdd/jH6icc20SMVFnqpPZDlziZ+8brS8LO/Wfh1jIypbAKuau46LEzHQHXjMxA6H/1XKiNB0yM
EhWpFgBE9I8HvbtlYBvxHfqObxxFW5egaGibm3QRGCdXgNrFgz9u/LZuuh4wEOl1kpUFimSP4CqY
Zt1g7UTzSAYxV0opSCYlf72ZwqWJtWzu07fBb7+Vua8+TUZwsip6lWceuVLdoPTVNGa/JjbByQLr
PL1wKrwcbPTAdaufAI9KDIaIv9cgRdJc8U4eh9bHIbih8/B9dP+yNUnTPd05ZRZxzhVXff2mnhwL
9qh4en9b2+qf4iyjx3RjaIekVTUcgtTOq5DdQddFQsvOxO77gmH5LYxwG7t1RVViSMx3BnXTAYIL
92Z6u33jqzuu/YgxN/msrKjpCObLclNE26tcA4b2gEM91euKw1c0pKbIeio2YB0L3nqy8nM8MDFz
MrYo3575UkNyH6fCTpugw5WhpOQ+d4rKVtgWSJ0HDUJ/FZSqcyiJKqGP7FBPWAeqS9EMhGS4/p0e
oo3drw9T5TltE6s9ab6VeG0PHvbl9sIZiljhQVNbGnHUCkn/YlA4BdnTecYonhjKElI7tLXYROM1
vD1IDos5QVswjwOHEf/9+hIa7WzFEtkgi5x3KimyjKpeHWuLU5ZClFr5bLh2OYqX17BJ1nduQon0
UUpg8iu36K14+htk65OITWPezCQoYaAI3hk3hV2sk398Pi8uADTihCQXKOumOfSvCAIOl7zl5agZ
sxDLU01dmnYJclSM4dapK6m4ykh0zElaQzvPg8xsLPsxoQtuju6s3y1O8Q6sQ1q2NQU+jacnXhM4
QkUgDWPE1lRgiBXu9OEwZzVMD4eseCv6RUmulSOOgU+UNO/zg69db1mHCkcTlpzvCpmMjrfcfyn5
QaaaBMAZi8ByJ56GKG8B4fNlKXI9LJXRYfsj77M+esFc8UeYXNNggoyJHgk3BPuu1hEM+Gu781PF
4keZYk89nNQLxq+Yu7Y+HeAI2JrkWXxr0eDg2ddzcO2LcZIuEDHSh+Istg2exnH3A6SD2FzQUQqY
uW7J3v0JAysB8cR3fiiVg7J4959JwljxU2xNKoVF2klMRXJMGkT8vk887hw5Q2suCS1ZRR6RqN+j
s7f13b0dYhjC6hom2Tl8RehPYPnM7P90pxHDa0YhwQ3Eqmhx0erPTuFiuMP+GwzYQH5gVBzUogQG
HO8CdZW3xhgxyl/3js22iHVzqSxCiIeLRL2IVu4tkKVVWJAp6AvN9iMvXtqAKM+zjHCGZlSS+uKt
PKyF/PuvwVjIpwhxWbC1pjbHZkQM2OQK9nMoTVxBDi3XuqxZdwkiBVa0Yr5K2vcqMdKuzpZCAqVw
LyyZkEZ/sIURkWs6M9u0D0qe/rzNT0sPbbijm82ykQXUxRFWarRBd5Ah4Ze7SQp91OFibK6vGUEd
M1lDGkNTGS+C7EAa9of32wKRFYEnwBuCqeodWhk3o6twXyfn+yWxdSVWIRdhilhLlbny+Wqv86CY
rmrWILQGe8eCghkSsWEjtXUsoDGwsKF4rnkF5uNMqNgjNvFtMG6vWaU2eEG53alvhxRAvpCRvBJB
0SWJz1tjueOfna9OuoDLyxNzU+DGbEEG7JFkEa+ilIMvBC9WtZcIwvGR4ON3RP20/2AYHOEQgwR1
fslQD9WHIJq5+mQu9+mM+Y+iVg+dkyd7sW/3pCvs85g8M+RC2+wMcavfMuyugrT0MNwVmEkXYIH7
hSxn6vM5VVAsqAiax43FgzKGM/YpPKdmsii1It6CTQa6T37rnF7WUbV0EMR9gIrV8ErAg9H60Je0
6N7KRAkjmWoaqdbdiLE//suL5TdmtxuEOSFDsb6Id3whUqflmwtarkLYC7tBsEKKgYhkfLmm1MBI
LrBL/SZMwnvaWqUUJN0rVtQFaBE3HPLHcqD1Qgd6ghPBN03CFFgN9yGMlwx4EQWvRuJkKih/wsUk
/NZvyJdvK+iGw7ubLCNYal/ATW24Ru9mVz4PGIE3KX2DxqOU1ZBhWRW/D1hKVrDcDNQrlW1GIzDf
Lsc4XcmWWJmcOhlgwDgFCzN+ij7EnBO6drGJREWrS1GgsLKjgaxO4JJAdR5kZ/XswgugE9pU9sBV
yjBYcyVcGZSZubrtGiL4Jw/6/p9r/VR7cCrCKviVocIdfBpSEwMTQTjvCZbMfPWm/rXs3FKZZYaZ
WC9Ohc+7Gvbn8qYC88Aw20UT3DvhEuneDJF6iLpDL2FuIux7eXzhegNEqHMc9Mrg9AJZq3w/FTSb
yJKrr3y8kYQoRqhXnzqn42elRgvsoLgs2O1SvPft85latfaN+TLgg0AnRo7pODD6VlqPdi2TK302
r1GryIbsftz1x+Uv9uN/cePiKUKuAs13wPy0viGsW2a8EukfLC04kD7Zuluyx0sAraiiFKuWe+oQ
juXSoC8gBK48CHdaQ4eZrt7DM1p91rWp27zEE+ZFVYP6v+VxmukSfe0KHEY/63LY7lvU/DYIzljG
TbZ/2fdVdKJsVLymPADjNaIKgXyv3NyVyqN7B089cQ3+Y10THsm5ssoZ7noXmZC7UWb+NFZfc4lu
gjX6kJEn8oqCkiOHoxiIAa7NeNelgIf98sLztZib/hfFzWkrQX876hDCtvRL3EySVB4RWHpSKOlr
+z83vxb9eRb+4SoR3UJvwIsFZ0gFYnpXZ0zatWld1Ck6y4gEQW+IG7Z6V3yrWamVambZLitLdxhN
6Eb58Qb/EzFA6l4tW1gM4a85/KhcpGSh+8cdBwA2L63+EgOgVCLn+KEBN9EkcQY3t4IoR3myvyMH
BefkoWrIgOgmvkZK+IMTqzcN5LfuVOoen8Qwt+61nNAmLCmpCa24K2omTM/XVC0sfxF0FXjBrT02
MbYPPXWnT8EboCmdcJVfz30O/fxHfeYM/p4t2QbkAPqraV3b228Sxt+6r4vt45SPdYyeLXoHY+PD
l1kvKlryV2/Dnsujehl4NrECoQ2uP3smq1y//WJNu+RUL2lTko2ypcOrQGtssFQ+NsViT+qn9fHp
BW2D3XPOt9gtW7ViW932wLonESeIdFqM9Z42KuyXgKUTjjImZCLjpm0R7p9v9GorNLc8GcCXTErN
12h8+eRkZG+iYVgaHVN4XGLvbMau/o8+Kj5+JqrXzKyH3L6gZSzRAVmB57H4p75oW4pXr2Bq7hqT
yshVw+gznGwmYvT587keVd3wv+Co/k91ZJg97eT61v9I+9LCskDfMA/mKsdm9wa5HNDn39nIzlGr
yBZY0ZQtF6GuVU0aVGy9gOM5oHK72OCv3TZd5RcZwerAmM+8SohVlHMLCrI+ShfS3XyicmbxxHGi
/9ddDfdyEBkoISUvHFaJBNGDwpwXiksjFF7USqMWROrzK1z+lJ30menmRV2H2fBPDS0pA0nX2+Mf
Bwdb5B2HUUyo2wKsjIFF6Hd3X3w8xuF3v2PGVeKeXiNxx4I+tH7bd0oLKkp7xKLkOuy7lA5e4AM4
wp6A6cQvk/HTFa/y5XsOxqjsUS8MyFQmGOBtUMceaC7Gqkg3m9ljYbpBiaMhTIFMivwQXbsXYZJg
dd8GGnI3fAy070ToVWhKzFFqHM7cKq6uaOFqdbnXqjxc3sDEd6tm6vQD4eYSHV8+IF6bKmxOwa5a
VdGicVHno9kZrzlmZIXkqFU30UOAOrepLpMrzZUWa//kZrRT7olQ8S3Ystz0CCTkzHhoCNDfMMlc
Z8XbbV9TBqkOmpIdfJSblFXX9M38D+/Rs1E+hIsHCRkePuU0vF1qFhpZ78tHF/38qfqqUaBvw6OQ
khQTRlouIQ0SoVcQH3xpTMhuOvyPS9SUmdOMl6xNSgxBS1fZXmz5oh3XjCphCpzgs7Z1VP/Ec6rK
CGy5fpgsCDCCBB6hvliaZQo0aRAlcV5stMzZWf7AA5lJmjvTHe6GjcDJMkJNQ4BrccF3uibat+vm
N2m6J7tzNdwkF+4Zx6PXUMcg1AQKkK/c6BUPGpdgoSkk2xvu92yfPOtUXi1gTq29usrRVCh9DKoz
Xw9e977CYf+iynXDhOpRwe7Mr5xuU9n+f+f8viwmF8RBn1FXHkyJgfqP97mR0NgxfuwHMHIFXmGO
4fOpFcTU16mtnykcZyWja9BJTvAgRwuMpAK8QAzjcvYXAVuiSUFM48lI1bkS2pECqz8ZEzgn3S5j
ZRtxlE2uvkIjyVt293YSTd3xj0/RJ4Xo3tbkucj/eG1S49K8vRYl93LeouUgmNn45S9bzI0HL0sN
z6hxEn/2Gj6JuEYWVZxG2/GkXzFgQktMAwGgHFW6BK1iuJodniv4C/r0yOXrCMd7SydDf4Qq9Zmp
XWctZQ0YOavyZ3wuiyNl+a0REBDkjAT03rZZ8TczCuzKzjNJoDI2Y31+yobzjnjUw6MPN3SV9cCl
lf++M5or8Htzw0B5pvmAiRHR6na+IIv1Ncou85j+tK/SK+K1aM79Pej05uRYAELiMHSh9FTJFvKW
t7NGfkR9IZko4c4wqXHT+kns2wtIJhxXEC8YLIzaj1F+YnDrjAMn21zea79p8bfHeaKsZtGz5teY
uACGFwtgO9h73aDTzEeUYh+IBXIITvkj+uXdJlVodA66bBhUJiFql8bH4gZpnXstfZYqlcV7nNmz
tSU5uXDuBoMs/Ho0FNcnJzOyDUnuy8HspWHyEKtj+ZN6jL1wrf2UuL7nNxhzgsaJMtcdmC7SWW/j
cN3dJh9cm6a830i8yudS8498SF5zgmR8HO1/QFTB24yVQiA9rL/xkvN2ElrBwp5P1Gg7T/X6W+5m
jFQC5w8E3XZC224GkGqllSWyC/HIA9yS/NL/ZVLXRdnI5AEs01lISdoU8i2JgV05CXQspvWUCXyN
qgG5KiMPTkGle/LG9VSQBmT6opqDoH63Wein5nuTZdp/S5/tqM97+Zo7uUwhdDdgzkfNpn88iwBH
Zyp/HvyU2v16I7ckz06jWAl5M+W4x8e2uVzyyiu3qdidwoXI2zyPpJ55FykFYJbjD9W/8RzpdI2B
KHgtaJ6Pj84dAXXXArR3wg27git30CPQCwA8entUz3ae7+Z5ZRjFLdxfD4+iHHYUf/UWoQOnpWEU
s7XjLOoOSrB9A6xYU1SpLUWJUr+q+kIB2n9fHOumDSQS93VQ0r1KOIy0zOMypd93Jr/3EPac0csY
X/BoCL3ij4K0cdYogSKOolhAKHtVnSZTpsr0Y7Je40PUJZembC8kq5VmwP935N/VqGnXk/GuTbD0
WpgV2GgEALjATmPQiKlvAol3wVs13JDqKlzcHzcKG2rAx2hqBOnXaKLpQ0V5t6BM/ej6zZIBrP+w
SuYto7u74GnV1lhp5I3L/Ou732d12vCx6FfjxgBi/QKEFFy43xSEdGhJ99cSL3DUD2CgxeWvKAFE
/4SryOfvAWYUj8i7rJBcBAUGIDKfvxwPPM5753t4m/rBNEtv5+qyvtnDpxhAs8rPXuGCAwXD8wO1
M8VglqUgwW/isp+5eGlAb1RH9/xnIFPPmfmAJYSVRpoGl6tQ9GuYTSwt1pcaQv40hTXtRfOTQeUr
MFfODiI3SOQWYWnrD82Kt9sd4DACyoZuhJhNJYCiWy0D3QOyehv9/x5MoZHod7t4aes2PkDn1WoB
jfkAIdOU0VoWwD39uxTzi8IkYTI1vVxQhgywy2T8xIDZo8Bm3qAicWXDFKJ2+RdzWXQQKNHRQsRh
TxmxdgoaYLIbPNIBX4cIpCZSi77V8SFiBDrhU37/YrEURbtgNeqMTLJAFLjnH3F+/fnq2nF4PaGE
Cd6yQ0EK/DZydVdTTW5JmiR0xsJ22NYmJiv7HhWHoBzNKEn/99ViNDYHyS65aNCZ9juSRCdapXA7
y+ABuzIxZs554MkpK94WFU/Zxo7ufrDSd8xxAhUULp9HhENI48iVysh7qSE1RqhC5bDopcZ2s7Ae
4Sayk2FV4mmffcYCp7TQmQy5rvp4rF+PHDWdhw+9GKKH6VrwS6cNmnzEJCxtgCx7Y4rJ5H1gnwzi
TzBuRWSeEWNajLWVGjpT/MdsX77yn7WHrt/2ZXtiPdP7rcnoRp3MTGn6BRhvz7Ligygs5qAWHHU4
rGbMd/T8+XkuXgoCIBeflKF7PYgiYXox7lRyXzghAyaJkH0Sgp4vsCyQmH9dPH4lpwy2JMVA+B0c
5f/2Kdqi4JgtlJC+YYApWP+q57veuoGlXNG8DRLTkmrJIkh5l+4ahiIGXTGEWhGFv8j6WcRKHVrU
dduc6FfZgkWn/6xuvuYyB6PTwDsLjP4D1pw+THMlQMbzsm0PSXCPv6/RGOTN/YkSFeIUEKm60E09
DlbmtujtnD4pwQtSZQE6PUPkyTU1HLxGDogErHOI2ML5o84RC8z1wR3DwmBstH6XAZ6EpJ4wAmwG
R+h/I09FOh/nMMSxWh8qlb3jJLkmE34TxZY1cqt62GjMTT6czgG64XLWl/sHtG4skh0lCUsViff3
n3oFuVJOh02mPHFBlLgNH6PAqQAQtYELzZcf8fyXWYXbJstw4OBd9UjSIjP6adN+GW0DOMLQd9II
yyJeQujQNH6SNBFN89bRXHq3qgDXuYZSqvXmckE0xLffxMmZCm4AsLhJidzEw5Hjk0BQM8VDoyJ+
wp4fJRZAuXGQ/Qix1zOBy1MkqrVu+9TC4fAU4wtnNY1ZxbGhNPA8u0a63q3mVZbrZCJawygFsqdT
dFBkdt/g7o7o34rRUHyUjmczT/Iz4yBAoZnKmFllNJ/Frah6iBCfeaCy/VOnMgZ/0NY3BVsepPFv
AF09eIqNzioVALvMRAhuR0fzEbPuKaA46AwKIZXl0Hw46jcRoiGj5Byd6UgSlBQZ2iW5hY6QrkkY
UJfon4t6wYtyNTu8Uq516WIjneaeeAS0AcYb4vkITtU99E0I++vT8zpUqvq1Oy3su7KvYqGFeTvh
Y21Gnhwsm0SWGfaAU2kc0nJTUU4MRVT1wqGfqs2IAGngQzg8AnwW4SRz4eFMtswjcYENCotnleUu
8y9w4vXE+0aN2arqifX6QJlKAdchdGM251SwtN+WWIxHFuVbw05yDoQwaFbus5G1Dpele7M47Smh
TTJEfxteL9e7TTphR8lovZNyCR8hJ5LFWjTLX5yKJoFOU0fJpvm7f7r+QWutMvFmA4rrD4fkNFa0
uo2jYMCAOZ3EQhCQ5Ol4V5qNTQvmf4ACHlwmh56YZKvmduaA4f0UmM4eDkZMTheDuA0MQ/PmaJIL
wuNPwBqjnn69H4eyYBQ2GBkd0HYEIcH9OWFmEL64TSlrqtNkhbVkwlVLzG8RdbdvoUG7BldnJtoL
02YVcSROwiSZcFDSLFv4Kz7y5FNJJ0zZ82YboZQaCa/dfgseX267Y8TmJdaD6VyK5+uwJUPFJD9a
Kpgfi7aNeeZwF4xNQxGWYVzTKM4XQgGG/pC6qi0I2w6i0oCpjLUtuvMKlpokv5j+uZRydD/6DRQp
GJwd1AvRdZ7jmuyanT/2LJ6PQq3IuSdbwLdUT9r1YTpL/E9ckeiesENxUmVgS4CQrAPlP9hNtheZ
2l8nJCi4wlWYgnxXT9lqHmbS/RJsFqAJWX1h7hhNGeQY4Y84ggjeQ4bml0HrXz0KfXKaJ7oTDTZ9
9ZQOeEiASAuxwoJv7s0p0fTOXjI41wrgf/UQn0jjOOjlxvVKfx+fA4eTj1MeYfoMUd+1/Y3zgP81
AY1WVNEgHaTC64AqSADIcwcUtef0hGrZPeaaedTt15BKXy71gkRxsUFwaj6KiplZx9vmFLmbUblB
PhqCROOIxjVdzJR3wBy63Ll/djFotA175CAAFwwOX7XeHSgx7JsP0Nz7GCkpfsthLA0DhPrRfG88
MexORIDCCchXOtZnsg2TpTF39EllFR0FvIU1IYx2eFEgfoV7VwQHufkVeIbwH9IX/BOCRVaMHyUs
dciHZxYBD+Ulnynrb8STrgre/S7/9FSTgsuzqzovuKcIwAxL0bsH1z7kByqSqaR5wnac9NK6mH2X
1ToFfwoFgzWZrbXjoT0+qKXm3W+2LU8/enrjEOOOwnTY095zsrcaf2S8ytWvLpbTe2d25dIwWZ7+
neY3tvoEFICNFC6gmTCcvoF7PNVNp/yn4DBSNghI6F3HCcvd8HrXNt6DKMu+cO4xaqtLs7ZbzR4c
DyFtE6tEdmP+J6Tvn600Bcg4nafjvctV7BHA6+ZIKoFsIGfiq5fK1uy/C2HhyG7hlsizpV0C8Qw1
luY2wNSJ4D4ndRxMu22WDD0OO8Uei6jpPE9wrkGssVO/mNhjwvwG36AtL4JAZdBBLdcJf8LSLZJd
pc05X0i1xsWS75nNlpiUlNesN3uF/UY8sEHtkwqwu8cYDV1Q11SKM8nEYXj0S7rZ/GIotXh9SYEW
9VZokSU5VyZ74r6uXU+h8AqYv81fQwoYA2Th44M2RYlnY0rqzRDTCiDOGIQHowmxSJ5UtitYkMzj
3+zVQojsHWOcskffdJqj071SsVuqvGuTvNybxnUVkSA9uqd/K6su93JKuFCjQSXq8vGV2O3R02Ap
06JtJWJcdZL2MvjR/DHYpYVSXBKtU+/xC9INucD3AiAZqMas5vw5GRD4EawEjMh2c0kbVbMOHqz7
qXdzwZX5RiaydCf4/guUqvAvaFvCzuGyDjcpUexFGOc5Bqt62S15fLYS/cLinFzMSo2NDQWzZnpp
h7XjTNkuurAjX3h3C7njxWwjLscSodWqFWUdD/QHZrV2SNkUu2SuBLvLbpsy3uOmXjV2N8D2qhaI
8AFG1AvEXh/RzTuKlzb5FUHz10TAuOE2ivbD6QCwlUqxrTjGfRUypytZ6wxbH3zp+1cpeCLnA4Ao
Ir0YmSAuWTSa+YVOzZCtM4LWzPXNRC04yuXJkqPJAigZMcjdst9VHaljSQz7EeyxJHVhNopH3+5f
+0G6Xx6TQHeW3csusalzNfJ2oxWz3J7maf+Xx/H9irI/Ctlsx6PxJUgVjgLHih6GRY5Q7aZJhK8+
yulP9h9tPgu5G4Y1zfy+1/iFwznFJZ5nZMKvN/EZSI1cuHON+ZOLBJMGocqQxUXn+//ddujSsj+I
8DU0dgXGVLqBCbLncpmNzjJHUkt1x7kIJ4U4mcSuTyjMU3T71XWPQ09ox3o0EozMxNLqMi6nlh9o
bHRKta7DuI8rrZ5A2RCJYH74J59ZoHqFwvUpa1AnZv13NfJEl+MDnhDwTqkV/0yCwpeJC8TxK3XO
aT86UqD1AJekFewzhzFMmLMdkKttoXE9Bql0KKKNrw4jaS2e9D4GyfofZY6MJCAkB7X30Oy0bjFS
XFnplf6XrpB6LuPmUWHYW0G1eSnEV58Ajpvaelb9ubNCQsZYwen+dXTfsLfZ0HpbbNPMam4r04SI
La32cLAWTQ418ki9PKy2OgGREeHFIODtX47ndLvNODnpctiArC05pTVy87slSkCW0j9sa+3kVB5s
HHAfQkFGWbQRU3qUzsjri7Pas6vEisHLgbLOrH244d75xnQwLYCEDJZyUQvB66ycxgcXq7qOAVY2
BG/hiRaOPHeq+bp3pdMoiUKwQWAJ85rG5N/0jV1u7DJ6bYvaRAbGUTrBf6JBwAixI4uawm+ZvE9M
gzS+7sUZLoeNsKbl+dS8QMKLrR5Q1xC7MhVaQlmUy91aCcnwxfrZLEKixYl5A9Uyi9Zob1ApNpyI
gYIu+UtiPrKzxtscJubNj1CAc5aPaRZgMuguyP9x4TQ5KAyzuETBFRtFdqFjnDQB0NLzhCktb6qR
trBmUIk5OjZl7XPt4Sv7v34pZggNM/56bYpLq/a4lLokrAcOsL1egimMmXbjVAZGH9N+Tw79hBz0
RipAfQypCP370WiN7pPqeWbncXi37oJ8m8yqj7wzbdFUDpxxqT3AxxUYdOMbPpWEttHYKsysgQ+9
X1XnMJchzHvAu5y6v6Y2/+mF9wnnmQ1M4N90TM4vwvdztGKiNAQHcgv5V6YZYyLQLf1jtAbyaImy
Gs9EtlEfwFdzRmhB86dGJm2rPd1rw/3pMJXKooqI5MsF0H6Z6gs351NDMyd4ICm4FQL1Hda7gJ9r
glR5aczqrT3boeo4P2S0vyaGIu0KEyjNg4NFMiAtIihoNSI/JCAx38qSpQXKRDBBqg63X+5d6hMQ
CtfZ3Ygmo+61iuG6qGzu9NQWIQVgGcQ222C+aN+IpAJ1K/feZ2bCs6BjH8yYWn40E0vV1KNdqyBd
upIkv/z+fkGFVGoqddMqi1og3I4yL7ijOR9WDAoYwOeCFg5usl32U9NMQ4sMGKwjPFoJAYVvgoOy
wCRXofTRK+7A5mX0rqWE8Oq5WaXXpqGtjlwCOfH7tR5MHxNawjgjq7eQzFXD8ge15f/h5ZpIcNWB
aKdDf4fyh8I0eLnmeHyKkeQu3cjnN6v32XhaTygjiNSDEGifHI2g60zNKwe9JfIW1GUvORk2cFAD
KVqNhvft3j+fEV4dAb03fgQSvZvipzmA85SlslfSFKfK+5FEIytHikAKgC8mssbzvX7Vem302KMa
637FWVZW740Xt5zQyiky/5ZFD2MmKxv7YXVSa1mvA9C3OXLXR6k9LErVv4cksJSWggcUssiGRzL/
VsvoNMeqoywtu01Qr6u0viZlL7yj1BVoXA5s9TghApUKC02CcctfVEIsqpAPzLKXs4Ska7fA3pdN
h6Aqy9PY49gk+2osO+2JQPsgnVQ3AoRwsN9bw/A+CMW3liPfU6DLnwwLhdKRhW6dBGv+YZmnxZh4
aoZsC9yGNYuT+ghnNXtTde7NC74UEzBGFf8QCSkUbMS6eS09NVcPibiP9UOj8sMLaV5oWeuoAQ3+
AB6K7negjI4woAORC7OMLpoEhWpm4AXiooK+iqEeQuHnjXuxeYILyJXnzx4TsGY6IybRcQQsFFzg
RGcpilmr90Av3kIKlCQ2sKgBJBOp5yqIGTntDR1BiJESf/TOBL+odnBiGaeGgY0idQbPlF+y3sgv
Y8jqGnbtoN7xSG7qQqYBnJvrnp3x4WQs+1JJSYccaPFVIUWcNR55BJtV4pH2znQXop70VHQ4+KCI
TWPRV9sZYkWUC90MTAC5xpIczr2TeYVwEvUQM5FppIHmo2fJh526496Lkf6OsG1wxF/GWbLOd7dV
BJ2NuSA+x2Klz2YUqXizDdoLOWNyr9Q6RcLTvaByKop9IVhmZySO/Efu87ecSg8hu2WMvfPSHFcs
/No+S3KlL9RYCraHA9punEYCHPb/z/ThVOC1SnUL7ILqYq7TLjxTd1UR61vwXYPWmSwliG9VZh2h
y2hh2XrUav9HpJ84NueYELrEKYbh1PQhOcnbDIRZZMjkhcK5+tM90ma9FW5VUNbUhiTI6/Xr+vzO
rk+8Y8uUoni2SXkzpJq3EYAayvqvxKiSXviZLNoQScF6InGBNlh5IWaJEbdBEoCNCXiVAAqB2YmT
t1VkH3Apgoj12zzA6naFSLNFHGx88yKXqEs14MY8lLzY0BK/uI8wN0NLKNFRZhBfUSreB080nqDt
Na9WGnCPM+85FWxaBxrYiFxQzkIDYRXlU7fvf8Yb3M5bfUoNnjKKQ7KN/jFXefLnuJtIlfEvVf4Z
BfNejO9kL4TscK8z/t2gYLm18ZKWqhp8nEsacy3lsFEnOyDB5srvR29C4GpQuDXy3WyXPET0EOZG
kwq5TdHJuCPd3pxtC7h7KrVmkFGicnh6X73ku3vrv2giinxm/kYkCvsfnw3kn9n0uaoszRnRidap
l12Ya7US4iRYUFib2omJL/dil2JgguiCUacIzG9cuinArFjCjUH7Q3BMj14Ocaq4VqsjebSUWP1T
1FkHitdyCeQ9mSLVM9pmHES6vckA+OFjDeF+32+WheGYUTB5e+FLmiklxRhnicjDsdBUNThugNAQ
2hyGyypZDwks5WNEcpyPhdTDLpthQU4p+2YaTOd1ObRgpNW+RsQ4YxwGp03FazLS/tUX6cqFUZ8w
VcwZ5s2ym90EWRvA9IxjkByYR1DoSkTuWH70FjDcCOJBSAmyMDurg4e9X+Cki2gcw9T3V9EXHKOg
EfvoVsxBhdOFBeX0Vq4FlFvGFajRv6FZwwDsUk7Eog90qhfbZ0zyPN+I9qVSDN9xo85vQKSLnRsq
DVET2uuZVhBwXu3mt8tpBx+4p29bc1XVddb3LlgEpdG868ohcvsNEifbX2Kt5Yu74CUY+Bu3cq0k
6TaLPWj8wgNUXXyuNlt6SbK9F1xWcDd5qdbQM3HLqhuJikcdW04I6Xbw2RVuu/AVX5CSFfCPTwB0
kNa0+pkj7GeQBohEw4to8Qnk64yZMPIqSRPBr7hBdLnAjv1/5rb6zrTVCOjn1EWcDWB/YTWQ8U8C
1S8rtPWHVqrJXY/EDeDdPFgg/F07x533bs79lTjp0dofuLp8/unDJgaVdJEA3htGxrMkejENNY1N
o+8CgQEaIXL5Nry9frIP3FyTSqsSK1xmU3hDHib3tN6kZ1Mrg1AjZrXV1Q9Q7nTqALqkjNikdI7H
AnaQY0gRismVWKq/hdPcWg/oARcKfCCEE1WZ1IvV8AzjtNB7la1jWDGvdhfLe2OPe1a2PVXVWBJB
wTIe/ktAhngnzpKOoWzJLVDcSfxdG5IeoaL5d/sI9FAFgVynx2gJ/Ivdj33Tb8HRhM4QYRSdpWk2
GyE5OkyD/g1Pm3A5wjJ57T8sKulg7Te0p94Xbs7/5xORktJIhIf6vwY9dsTic4mj8X8uJEPI3S26
UpFN9sQP8wCm+9wAFNwWvqNTNBAg+yJnzRooZVVqIMX1TGbSFDjRahUrcIQ4+ewDi9QJPWizGFTp
Y2/V9MqzWcwULV6u4yvx6qLe923xlyGjCS86/ATuRcFFkDdAtqAaYA70HySBll7d00JDvoaaz+Z7
MYqJyQu7JSGDocbW3Lk+kgCgBRHEQZOfk7Tk9Ord6uOtpPcRgtjnKBRpCKw/ibQ4i6it0SHH/Wlx
G+ddC9+rIZzVbNMLgu1e6Ec1FEQ+LCzUJPZIruOZiBwgk53CPwsOfBJt8A/ZTi5EDvc+Z2apGQzK
Fry4e7VS7wO7lYUerxROruQkmL1Bq5R4AFHviAuzvRVEIwII5TL91XRwT1qRXByKYNvZ8+TTLDO8
APefCeYJ7cvtBG29C7/vuDCcdDMpVc2491muAl2mRN4cXvuMi/6mwvZZvD/SJAyhK1vrbxsJcWbO
JrWsbvbUoQJ+jjhQxxe2xgbNqYbdMWivslGQ/wwlVjBam5Os0vLRPR3mU8lSiPqylJDqV7vBx2Ko
13q/LnxWQ9Ghl7Xc0uVak7fpqOERqqcyY6uF3Nu3xBcHXKWufX5zdJwS/X7vTAp1OSW6ix0DRls2
Gp9jw5QTGJQOs7Qhidg6rpMb2HNJ6XcNY3VE1DJhoz4dtol6220fW1KxezAO42/GVQ1TBbtxCS/y
xUH4F3DkHYcOE20Z0I19nLAij6j40qmx+lRKPwx9FzIQE2bziifxYDNwgg6oiWsCpVk7DQuQGeFA
+SKT8+SAabxpqwwgSul6FQtAKSWLIjs7DzO99iy88pOZ/EMPXEI2SQ1vki0RZ8VYPqKXUMdgXDFp
6/gVdUMhoFlt5a3MXtohR7LiLseD0/Np1Mg32GRjH8KilfH2QtlhUcatur+3csET0UJ33i0G14hg
Tmp3MFgT299zi09sFepM7GgxnX+jQo17Ni14TLcgXl07/ZSQg8suloEkJxbApu5tzzLbr4dlRdSl
M7uPwVW19kmMRmElxwdywOgMFo/ztn0ajfFsmd8AjrYdCNTOPX/psHtrb1NcfAkrB2QhcAW6gvY4
BX2R0Bbiwz0sgn+Ik34sya2BYWzg2JCivRctJbS2PXRbuV4f28e0toObX5HBLWnrsDt7itWzFJFC
gL74HOd8Da6BEqYW3NVAagm1TlzO/oykKbBD1pBvoufj7eDQlElMJfet0AZnZQL4c4YGyv0RGn6/
h5wfugL1HvsXAux7g4fY0rNomcTwCOyh/s+gJnHmVimcYqanMQKOwk+bKcGYDf5ShUAJK6NVdC7d
dgT+h4KN72n7BsHyy4RmxXhkt41w7rZYWTp5EzgXKQAUN0p8ddM0sE260WrKhuZQU6puQZCDcbsf
iaqvG5buBsOsbccK3IorbDJtLtTw64j1NFYw2r1eqGcTZxwGQQsyw9xpnWLr1fuXPiyZ7Lr3lWoM
Mm2FJwOhoo7Ko+KK+UhBWowIZUuLNSERXmV55UjJTbUAmPtv5K9KhyEzFs7XIBR4A+dP5/MTVak2
thdIs5nC6xWWIh7brPKKzqyvvFxkz5FadCcWr6nbgtASg74pRvCz6brvfjxMoWjUBdERwlm1OXKl
977kBUFj8ryo9DwB00Q5Hkb8zgBtkNQgr60YQD00TTVk01hXw5qVwP84Edr4Rhs9o58I0J9f0F/b
br0UcorKszynBCbKqorNQfolUPxDdN3c7nfe+m/jcBn7Zo6SkozhqFrv3JdvJ+N4N0esE7Rlfxm0
r/NVRYbENfkxxPq5gyCbi2wJV0vRlHKD226pSbsR+6daudeeYDZrgabRz1D0pkLvo71xRJ9Iia00
gvCxFdz+Va0ci/rQia2pBbXtbJ6BRmfjlp7zCQRGYrGr4oob3yPtCIxqKHoSucPytz18aAqKGCvh
2KXyGfR9I4zTouiamB1IPir2uYJzgPcvPji7NdjYHRerJMFSShtXq6p0BiOq8i6CSyFJsefe14oZ
+4Z2ICJB7Vas/Q4BVHC6YeSnzfSuRVK6B3gZj64nE0dOFFecrvS9bjxRatgNwkFSds28QxkUfqZ0
R3GwnIAeiRUY+15bhxI8r976M+OFioe+dZ4dXzISqHrlSQIPo+MdF6oVKsokDUa0nmpubL13Woh6
9h+FRBGowqXhUl/cgAbpzl4zvhqkmTdU6q36XJcm7eGdy1nUc8CQOF9aYhpdXS5JCYng0Ws2mITR
HMws9TQJ62aSfJ3Q0ss3PD3HnKSSRrc3r91S02DtnyGxzsEMYvtFDZDjBwiLgTArAKzZGygiB7Lj
i5ZTRiFgFs5PkV2CDMlgPKwhh7lBxt0EM+R4ENk1Q7/7SoTirYOZpKsxC88EY7Y/wwVSoC12aKQe
iiPjA0eqZU1YAW+FFCJtmzcyilkqXNCNepXEvnz9ETkIxnXTtxIbM0rDPwgfyncFU6VJZdeAC2b2
y3wEEkvBk39SgYKziLsCpTwwnr1DLPdTZ3LM3Enenk88N226ip8GOHZ4QTzakq15SGcV01h+U4Zo
QlIgfFsteygtCnoRj/hWJpUUW+bicTcpFc6hFuDaWdnv6wGNxj1ZJUtAuUYpEnDG8Ckzy4qnkaWp
WlLYYFcJzSK/lR/LUqHUaslmWGPYcQgeSUQ2nmNKQZISpN7ZMsWx7uIBABf5M0XX7hfeClzOfxUq
ipZqvuhwoqmyidIH/bZglU4+qWhckbAdVwUWtXq8WE+XTgyE3U3x/Qh4Li319Y1XKzOa+qgUmOrM
WAvaaTlDUwnvlB2PKnobRrMk/ydZh9oDPITFfLdFqUOACYthYZhPV4GqMV7jkW2QgNCXj16p1Fm0
EaZ1il/mNhqeoGU77T6hdW0LJV0QVZALOv9knQe2PcOQ4y6NEcTvpXR0fPN5slj4Hesr8WFczlAX
WH5J8xev4o4z6POlvxT8rSc8C2ZEkgRdbE15bcYNqeqCkImwQ04Ew9xq9KTxgcLdVhpx73tGn2Yz
HNfp1/ZsD8k1XiyXBWQ3xxztv8LkUBJXFgpaW23eW6WcheFs4bvR+UuxD+wFSy1VsuZt3bo3nDcG
jpLOavZmLRSGtvx7EeMqrrHWBymmLS5jsbZYhhfKc6Xq55TSyQf4dwK1qY90L0SEu/QzGp9e/n08
cPdWMARnnf/LhutCh0BB//EdkiGOsdwFegAun1Yul8p4s5gyOEahm6eXGO+LEjtPufm6IH3NX2n3
G7/c6urkAWJ9xkiiGxcC1tWByCac9e+JI+3av8oYBe3mUK1duYjG56jWgAnco0sELed1pV1N6y6B
BZTAm1trgsUi6u9jQycoBj0JTGJCjflQyKUoS4B/SijmRbZW7bOSkOO+sb8WfS+NEdlewGDQi9Nq
CGPWL2/PtoN6xGXULmSveVK+gdlerdzoNFO9oLn77axK5Q4K4ucRCA2ifV46c5jL54ALEVCYiYXS
ADHvXM6QQfkGZDrgddpL5cn42K4soZpK61CkeGdGRD1MZSxp/KHM8Hhdk+ni72CshTgXNVQp36B7
dRuviq7D1P0i1+nB66PDEB5bobx+J7G2QxcvpnQ8us58pMPRG5CKHzwk0o0WkToWU9PsX3ASikzn
Pz6zdVEB2QNrgFP2Wtr6sj31prPZmduTpJDiRmk4vMzC8OqqTkUT9YBDX6/hlvbHoaIUIa619AzW
c8HkxyV5u/jjzkgzv3XEd608MZYdhWudf3zM8O+ub/Fpig/CYZg2Ah6ldZWG3OzG0/q/XVajGkcZ
d3bApp6z5AYxBtWdW1MS0XVaPKkODshH00Ek43OY8tXLZ7u3FaoPV4F2B/I/COMY3h9NtbfL7zUt
+IQAm5dGAl2x03yykpxd6incTT2+gi++1NVla6L3Hzz/usF7OrPsopGWKj808lvqeLD1p3k1AdTL
2Lde4UT/RyAi6We4GuYc+7x9uSUCel7i3F8ogE4cBmZ599pB5ol0WxtWfy4aGLNSUNN3d4zxpoX1
GRqFXdOgBp9G8J2YvEUqor68QBbK73qkgGxLMJrMCuvNAvO2QlspRPY/yEhXtacb6/wvPens5XcK
h9VvGWbefg+82AXooBDQsDbZWFL+OvwmmlkXbO0ydjj6lHfYqoSYt6k57+UeSF3RLz3GlOpBUCgO
mMRg/8i6C52wjahQ/9ORF2ybQWWdP25W4ZOjubF9YYFjD5Nvz1sV1EJB1mir6Jc9A8unYInyU/YC
z3KAWaBswrni44mxxCBjSTtnx3jtM7meC1+pVJjaOTEFauwXcMUO8eUUIiNfNPNnqzg7JjAVzupK
FMfN4XX7n6pUtXH2vB6LZK82qbJVkiE/ELdUG/ViEUciH2SlRBsMRovSjzjkpleRQnF4K56c1dyN
XceXF9X5v6HWG1+bepSDnrPCMCOZT9l7hDT/xub0aKObJG38FkV6993Q7OHD/9DoT40uNDDAL6Pq
WQq7P55Uttii7nksn+bg3GDFDX+EMAuSG6jswzqSv6aVgS5pAB4cXZko7rTUXyhDGXPdHTv1UdKP
63ibiUH3+Xj3Pfd40axPxUk055ZWTrfKr9DtAwN3S4k2RhjeZ+bDfy//d4U9cvyzOLnpV/DuM+E7
I8y75oMCeR1lsvzsWD0bWieSCHOLr+HH9iyi7W+uGopZvunK1ZkZFOQz+g2kmDZNtRP1SHJiyo8x
6aC2hoiVNP5ZjqTx209dushrHBXhunO6+yPDafbawjTkB9t4fsVkh1r1y/134y48ayJNbGRNwccm
bXMq+NP6+eMkYAaP2LYpoze3MBKmzsJpAB/CkAbGuXi9YDFI1QZPUCwrqgj89NOjHQRw9j2lc8RR
cvX4OZfvqKIMcmvAnA2yBNWSTjyNewZntLqM9moHcJXlkwQ+fUq5GGeXMEN3GtT8S9hhFma0BST9
Rd3uChN4RqtlbT/1L4YNP6fPutz1otY3qBiN5XsW1faoe6RXKfORCiV5SaIRgXxDyW3LZe4j5y0h
d4nUA1+fgPZqmCRUEGDavXNgdhDy26HKdCbdrcReIKpZYmPhVC7hbkgShEV6wGAlRKFj9BLLcxyu
X3IO92Ahkn44oH6PIGqE2GGletLsg4ipb6Zq8qP7unxpvOUjRin7OhOjt77sPgI+wd7ewEWBFnvM
HAqZHXyOCCoG4RCtsIysQnRB5Ho6l7lg72WJ6lpjsrnhDUoaIA8po0d/Y/KK57jd4weNpjsQJdgx
RYWlzdoOAjHlyn3A+QMA5BB/Vqr6L6jYhw1wbnoapULYwcMLO5WvvAg5NoYzfWQmJrd3SqU60c6s
FRvXEjZB5O8sAIw/0QMxYBa5OvUCJplh/rIXNzPsvpDWwNrvltfofbarsv0QZIYkZI5VQwhxwk7p
JgrV1fo+G23usqRxe127J4uItI3ba22zOp9CcYee6bDTzo43MFHScF5G0QSnynwwTh9D0N/sCs5l
eRPnwjBIV72gY768SAmP7bacY0+VtBh0vJY0wKpLsDzTRdzqFEl5r+rKTchgbBQPj6cTnB5FBaHR
1hwDJp9wbbbrzsAsg1i1gDkBjiWVKqOP3GQc4UgxpwDrE5M29VfTOSm96U02UgaR0ZeAVGsE2hnQ
sCivIVZfEpg8XmtK2+cnfVc07g9LTl/gIT0tqZ9L+6YvMo4bVSMXcUdu7Z7kQLaZWizmWV/O5Gl1
3wTL+RExnbB6x4P/NfT++v8Axkv87ojG6ZwEQIvsoXdotG8O3MZOCML/wPeLOLoUQCewBtL48dO6
fbFV3LxR/85615GIdkf4gyLJymqnn8WYTy6Gp80KhwCrEyqQ0UifpFou2bJBEG0hIHowtauwKHKN
wllMNPKV9Lv9llRLJ3y15UuvWpXuVRkFPtb9GqkC/xIYEH5TTUOB3jlodNEfC2Gh2zTgjlUKhA3s
EhEN9NN91FfmzzqsOzOjgY0zF3r7NrzjyuTVH4weUECTMEi/+s4PAtbXZdIhet/VDWxODVsyYJr3
mOVTVtOOYdGftfEMDZBPzK7ES3rs+Loh1gLL0gp25sZkyh0/YI5VNSq6DJLupVFhddTlq39Ch14s
w3629spYtF2SbbTq1dR4SIJzeNAUVYI9Ab+cNx1B21JqooLdOXQbOdf7q9ghG22g5dpyGOmxki7d
7sanF5PzDIXkDl/DEutyEy6C8BvZPDQE+pwwxl90rNLq1wKFa9upx4fo7iYZiQHHh/tYhwF+6cCY
rEIWwIVIZunFtKIKaVsO+iStLKHdoXeeSWt83FtbzUy7JHHUJA4Ake+N9G6rKfFyto/BPPT4ZN7t
KDU0ogo868D1Rd1gdj2lus6/0b4hpNpPUUZ13i5c1dEhpcNBnMOIkywDhePNMptbU2/idKkesLFi
HldxMtMKiGWiP13p1OWFrLPPvH0vJDv+LD4+luRd6e2fVvQ6mKmbQFwJvYQymrXt19jj9y2GqGBG
fynagE5oR/EVhuXTlRMrvb+md2l4yp/hT8wUXLCjLdPrpto6gnJwUP6pXSlvx9R+kW4DLsraA1bQ
+h+K3jNvFDbGWpFfvE6O17BPof1/I7hXF+lINqNZ+6s3f2Rl2DR0uH00CWyZ4tXJTnXsywrD5EUl
6Q4Q0LKfwI6U8abedOLw/35qkhJBqNprBCO+c+JPYJbk6XBK8GPQOvXccQKxfx9R9e5d7PvneRbT
QlIiH02HMwf5idtkP6Va8TNuai7E5Z++xarQ2EC/KynZcWlJl6lYJHqJraajsMfOWQcsmi8I12Es
ycz2KdT5Eb2/NaIT9vQpFG8Vyv2Z7XRHR2LFbgvShJhRq8ZY7Ap7w8lhdRC+so1ubdnjNzuhZ0RJ
LtGcRvyLH2ZqNRAj+EilFTnslbuQ45gDTz1wtVLy+OFe1m/JxQo3/oF28yibp4qubVDRVXvcNSgd
KN6DkWGRtaGhGL6uHcuXeJ4qDBYRrfl2QJbTnFA+FcT4lmXY3ienotMvmwVzfn1IQ/oPI55fMUyf
u2MzMyzTXkHbp2MAsjsdlruvvryLo2TAFO1elaRX8mIkjM0BcQi2al1LjePUhxRpLvIlAsuXqCA+
+PYHyISiuga+1nDfYmIMg/5e7hafLnrdokl+3HocZTkU6EDMc/Yl4yT9p59MErT4EEcYTn35pMse
WH8fFsKkz+jlC90SRKyndvD9iUOK+EQvWmJCx8wsBRwhRBkIrN4RXlaMSvfBqiz4CA1iqfrzGTb8
qXYTxAXIf5kFMMjUjunHGiARKA+KUnM1bIvnw32B93VqtiJMh2lWGQwMeIpO3f19kXoUCf3JczKZ
o/Q5rUm5sCKOyY7wxFKZjGC3EduCTYfyCUAWExTkLkWd3HFV+6HIp6KYWdAHHpPubUJD0fWrA0ki
QsheTBXNqUVBtloGFQSmY6F8mnw8cdLBWeL8dAeGj+zcoa8I0InGKow6asFNQyATpy/expp+Xps7
ybruiTrslFVasKljn467Bhf6efKAroEfACvHUysNcKsqWiSWt+OJaI/i3aAS24oaAZYoJXabaeWn
1cgV1qiEh51LcuelPg1feyL6kAkKM6OrstPFVrLdmlbHiXEebJs9DFpfJjAnqQt1d2zWLxTllN6N
r/T6bnJkf5q/yAWM5567s8JgGeuZCCwB7nJ2BdWHyIRF1MkHXW0hCXIcLAjIoiLPvE/nKB1C9Lzr
6222W8cO9cYufEtnQ/dYf8dvKRqF6ZRJIn+Vlmn6NaKsTBCP11D2a54H4/76jNQzP/VKSbcuersH
VY5zixD98xTgFeDTPL2BHSNF2TLNU7PIxqZLrW96kcyl9N/tPA2/ov79xwsi/xPcKXcBfS4d+sGP
7Cqr0qEzvxxB9cBZQeAqjv62uLl5+m2YRxdLInHP6XFvfuM8dv3GO82Q7lmWxKdG+byTcdjKhrri
vTU7bQkUt2W+wcRXPQNb1ulLqW1XDhEZUYWX3hVk4rMH7Jrn9KxbW6oo/lqqDjG69ZfGPOsj8piM
qv8hzWXee6vuck9PYdwQK5+8dw6PPH5jiloFTqQqVNlr38wQHm3/zfc/ZBCcyCrEGLLg3p6ua423
WyGA2bPHAxJ4xj8X2W9R7uyasnuj7mj/O6sDvY1ySkqwzaSd6fD5hNIFVl9VdiwoJwXzTGS7LiqP
pcMlgD9gup1YUGa4Hpszg53qQrKSkojbqTID4VcuMq4T/SeqOsX9pNrQ0ReCWf9B9wj/ur2QFh7T
Bt3IpwGXRHuvJXR+zj8KkmRmdi5YjwroHT+fv+Zhjp3x55i97jCZEbiwwBATBrquao923tOP4AQq
9VxbMFeaKamkZl2u5IJbzf6xIw0wyvUbSe/SZAd9zS9mShG/fGrNkN6QdpM9+5BbtBK1muGY4YAo
HIPz05QmWu2EAC86U6TbgPfDpxLJ3q1C/MtV4IfOotfmGaRRae8oKkpaQzfuzZRgTTObYpl9Ffy6
YZuylJn6DdPiVEH2JDFma74crg6TwDk+BpxpZjovFWpR+XjSYdj2oDqH61i05ZXVKRJU99kmd3N+
bfH/ioKh5Q4QTQWuvQ8WR8WssZqMnD44R1/en/ppy/Jnh5TAmhSNM/4nRbIMpDHaoxrkpKi8WYWF
6yd7DgDvsFsmy3a89PJF/8666s9JoIQay/O9BE9zgc1V9es7l4duAz/yrgQr6xu4GjCsgeEHg/E8
fuCcGf8xDDMT5Ans+Ha8XTTyLF4jWSDttGdXBGKJErAYJ37YRnA159gf791sYA6Y2jTXOXSeI1XN
GKjx0njb4GFOwo9qTY7TEsTrxEy5OOB3SBKlG2aT15clWwOGYSHQ5Pmo/odsYpfzWeV78sMf2CO2
tcDCJwos1tn09D00ZCbUpwubi6YXbVBY/+edFHWc3g6jO7ytcwIid23F+vJ27V4X6yZXIeQfHmBM
WTEg8NwvPzPOzzYsfahO46oIu+esMzU00C5550icoqQE+dnNSCnz8RN1Ny29zaGRis6cdGfQzeBt
u2wBOIVlsCyGyy41MBvxfHFUureEy9RcPssUewQmEfwE/2NdEoYS/h7PfIdqdDh3cs3KnMtifHPJ
eOLtCVSR2IMdWatk5EILjav8IN5a9caSwXBnV2eB8QsbblLx51eM2j27Uipx2726ISNAD1nAtzwJ
UnQTOgBLCCQTyUph4HKzLUlK9ylnf0/wuSJFpRQJb4YIUxPQ4F8WoR/93WzVhUHeowiR79Szg0Bs
KGOyWxKiCtKK40S7xtQlhsiB+g9F0YrM8z0P+AyuHAH7tgb8Jrnrukpr3SrDoOsd+0aXDWh+8SlL
lXQ54/sPZMHabctrQH+yq7TKXmJ+6J2TfZbiwlwGMFDC8W2UT5bxg5omYcWrV2Q25+8Prl3VQrfc
RUEiT8oK6060PXk6KkBOWKpySaD2AEhTCH4YLaR1a8VCT3z4CB6TKtz05g7CaQFgpz7XyB6br2WO
BWIfy28vWABV9/bUhKrqvx4WhGwcPK+eFcNB132I0udzz/y6ljYNkU6bpSl7mNQGFBIEchUb5Cna
xChcfOCDP6+xbsH5LwNqajqXG5j+/v23kPfY3Co5xyjJABJY5Bc81auiPZPlQG1BgTSzobLRpZ0l
I2XekQ7C/f1cL2Nb43ZGNERsBVI8HEU993rNQ1kM5yft3Dnbv6qClMKOe7xmCtGz45bzAdE1RmCk
LPnHO+9lioPbPVaSI3KCYFfHMDFx6ebJuPWKulVl1lWg8ggUUnpE3stC/Rm9wYZBtohHmzoY9ljy
eE4ClJCXEq8q5BU3YW7r7qoxu97ukOUMBtaDIPtO1SUT7Nu1TMHyGSKPVRNVPvdZMfW4R5eg245z
H2JI9t0kQ/09pNitSfEyYHjs4zGgjwH9gnSaqRm1nvJI0VJ9dyTdWjTAYew+Lch6uFjuIv5sXJr8
8x+SM7377uqGEj4l2DGqZRVcr2epri0NvXVV5xu4lwUarmRAss79fKdJRDvyo65iOkIG/7ASO9Dm
86OZv+adgFPnMz5U7X5HEQGwnD0DbA/2/UztFJ39800YG8DhHnyO0whLk+La0varVa8BlY/bmbiU
TPTfAZ7OOAVGbZ+h2Ea19Eepf6Bf20T/aEnR24P/OxRfqZAV1pUm7d34pxq3yhalY2ILYSm/bJDP
1Vkt6ZDTIYPRRlz7I6DpRHm59N42EnWKpyN7CK7iuS5/v9hVc7fBi/ZCtzfNdqGrOVjfsJDy1b44
SxjF32tZ/8ExqKURFhM8/UHMyZAgI7jnKL2itfUOXN0zSs3fKQJ6add1lV/NIv/eD16xT0y2EMtb
LbTmC8SjEJ/H1nlqVsbAlOVEaAp2t+Y6YJ3TWXLxKNXt0UNBeD6iGXPITMdPpC5hcMxtSsqa6lCl
7DyUBcPPcH4zl6PYIxHfaK8kGlzJzB21GqIgh+wqkAZg6QETNHH4ByZZ+rOyTvTUbNjOMy+Ej214
UrBhq7b7sQO6NAkAuakm2K1TMSzDLZw01FppliYLccqxtjcd+v4mAsNPoR7mo5ktLsU5MOlERW2n
1P+WDDhN8gocl6HSWlNqgpFzY0q1R2LejeWlqj9/I/8fUKk5mYCwssBeGxedVsKdQ5pIA4sGRzFJ
N8ze7QOk7bygwjZBTLcTmJL9sbzizgyPIhY1H7bn1b8r0lPfUk2v8RF1Icwe1+KXcgfleNVtt8lF
QzMMIamnTfr5tNdpcsz5jI1VFd5SRjBk4SrltOxYiohGSKt/YygrjipEC2IUQePuMYXSmENknFUk
vbXsU6rZdNmvQ0gxnY5Aq/CFJvoBOTZ50KCbRjylk4uxbdu1+/xMWhuCJZNsNlp6Q9M6Dr06se8T
1DqqFl4Sm7NPLor+9bDV82rFVVPaoyZwqxAqMKjhpAtmL/eo3MXHEP71Muo8+pkMIFiqTI7gbd7H
91GJBC0fzDdJOEAiqsHSb2RlkaxapBFySl3Arsinui95oYVNA3HzcF+BVP2o/GMSd+d0jkdM8k3r
wL1AAlI4a8hsl8vgLDb4jcSohaxEMz5F9TWU175WpC8Qm6fxDIh50Txr2dG2URTCT4VvjlCQt2/v
IAz4GOX5YhOaNv6IRW4BiPkp7ONWD79vD9iyCOPrDHaONZDVQdFfxUvyLg/33+UUXc1cxtH8vG3i
BQnCYPn67YroobBPzQ1ZXi5s20zmmSwPffrVY1K+nxh4A7noSJZ0uNJmMrAQDUAliCYk3e4fykFP
5AFjzVmu1AlughvarcXO27nM27tvoeOKGES8rOZpUjX7pEBof2E37XLOgx2yUVR2yPu83VDeLXMw
AzM/mm3H3KRwnXImFOaehft18pyWd8/XwxpQ1HU2mssOo2FcWqp+3X3IHMLu45vkce7GYuepTtZV
bBKDuR/eJttiz0PzoWAvCfp98GzBbnDwmNv7gf3JZ7v7Q5/7xBgoT1qnisQzJx5pmyhYmTob4BTh
+9wof3cC86cU2IvdnhmVLCropWd3oZ/odOVqaiCI2eUwJp01EEUL5BjB8zYc+5GyT3UbtXR2hUTC
1D6dfcQifUOpMFWi3Sy+2JUH/dWjuEkxDti3De4tbu2bcjsQ7BGYvyaz09h0mHDGPX0DebjLQuop
WQHHEG3qfom6xk0mJ5w9qFqVgbuM4t23/BIROL8KcyLyJ/jR5aPFsoYfLbDeOoMFBqYxuD8u6GF+
/73EHtlcnP2v8f4WbfUVxZJrS/uxopon4jQwMIgqQO1an+kqIcFxRhyvN7CWJGKi7sWf/9Hwlrrx
rlEgObgxUPCB0xuZNvyBBq3sreGtuVKfLWDw+dAFy7K+t0Rqt+Wh+INo4RP+Umn4axBEs/l3l5Sl
xJTvvbeK4s7xDtddlBWd8Vukmih63IYeXxRPW91UQrXZcYoT93mB+Z1hawi7Odp4R0KH/1cG06J7
ABoYiHwgVxAvjWYCgQOj0FII6r6+36qXwsvI1x+ojr2Zdl3Eb9ross6BfMdd4DqSRMF6ZeAsDihl
QQkdS4zgR0hY0c6QTA6cfsl6VCvyGjySv4413OGwR3Je43e/s58FnALfFHT0M68B2nmbtAhUxzTE
CciBLuEkOoqaWMQo/Tdom7rm7k31rAo2mVCYgQyD2rSkrA3rszNRJu8P//Mns+Ah2SN5TgUqCyt9
f5ncyOJHP+NzYegUe9/7FxJv9Uwu0bNfrwGuWKD4mQC9kszmMu6QPd7ae8J5t0/GTJ3hof6JEUrJ
4e4ZSfVSmtzXaDvOQ1K9nmitVBhFaOfEBpTSn5fHwoqjcVWv8i1tMFTEQreLwAilyVf3cmrQPQ3q
23KAgQYof9ku775su+1w0+G2JnuIkznoDIpvky3UWUogfC1ro1hFhJ44300XjhQkGFEAsr1QAIxJ
kJ3QcYcrmmhgo+bt+Nz3+qps4WXbZncJEBUul3LXmqXTgM6lOOxYJmd+e6oO+Wkhwde5Vej4m86P
f7rmb0bXrVD54ogAUxQyHlTVw4tQsxaCwHcW+xymYQjASfNS5R1bXgtxh13cjUdoNYQNg+g3Q3qP
GPw8e+lB8g8GFmf6ix4blx9oDx2bAWt5paIfKWTJFK23ZpVwqA7eBAb+uqEoKwGiSfa4+O2UAdZ4
geS9tSf5qhkCo0asYzZCIvXrwjpWWgtOeM6jNNdFcvZEpPWegW/YWaPkXusm8UJwhhp+P+fTfmhe
4KIV3x8iimVgF8FflZZXB30QYmbWz94RutACi8vqra2UpVzkOZG9Wgb+oJXvNL6o4gouh07G1G3C
viGRE+qF0z3pJl0gFmsxPImAFV5yeoxJKR8vJ0YclyRy8f2uyIE3YLohsqnr/Kle1KQ/Z8Y99wUS
mOo6VhSv2uCef/kMfERKYY02mHvBgEL7LUKymoGh+2dKE+hpdg+OSrek1e/fO4UbrJO10upBSgtq
rpubyxZECGFpmn5hDwJek70idff7PAsjyKprwdW1dqyrXIjzVat1KrD+h3ffAulTec7dK3Ig7Sfv
xzjm4tLLAIHxwQimTWqhd2VXsiLSKLmZqCns5bMqPPp/FzfiIcwcz6DSRQO/kB6Ulg64gPTEfXUz
z1BrQnsNMPTQsc9aTuwowYoTx5jedmL2AwByvNTHcXEmWDfD5onRWv869siS0cTvCtwRlGf1ETDQ
tOVa22O0QHNLIHpkurwl7SStAEjPfcv6fTGRkk0yl4TgGFRFXrFUvGoTwNB2fwKDQb3GVPcZax1+
V8VSOz5AuxhKD3OlbGXUDHWBeHOUugZ4tvs4pCZ+n2SWyKBqz5I0Qug8XQKRtay7iAQrXoE3+b9F
rIH4ZeBUt+PTbTP1DtbHeZITMts53yDzt5jf7askNJvTcKvtnzaDgRunQS4Hx1Ye6wpFBsGTVkBH
oDpxqOfEEYx18Kuge4xeOhana0847x0DcX80o/VhX7AsN5YMkbcktRsV01HyDgdB8tkwUt/l9hyl
Wv9QOXxC5LPhcGm0ZjDT6OwZq2PIRFPzokMWx1k+45edMet9h8PhTOGwrBhlArXuWv0CGlODFXHG
w74kvjqtGTfCNIlgMG144eJnE85tvt3maWMTpOSKqHg5DooD5uohnacubUynOw8PyF3swrXdwTpp
MvvOxaGna5yIsoqVHf7m9Z7ooVdn3Gdn/6N66PKXDHyZixBWUjISMNqjXZSV1SVfUzOSvQAUcI0t
uuzTrTAcuJtA5ZGrlPsYLV45P3KXD4nJLm5AXQfnEFeNHoRi0WmapdtUzNsBpIj8IfxYcW7FH94X
/dLrYuFnYx4OBEaJ/h3xWFX6HJ6TbvpU9WkiTHC1yX0cHfBH4kqlDNN492sVuJSHuyB7MkJJK9zL
5EpJXK4BmJ23H7fehx9qXOQmbiv5kOi8VbDOuIhJcB5XXbgNtjFh47NSIQ4OC39QAmzJtg67QcVd
G8ecx1BlBmV0q1ORizogM92ko+e7ESqhJhYoBqtoNdE1fwcdOCvlt2TBcMTIUDO+XDbC/0sNEg8H
rlUh2N19kJf0V+rqmZBvNnVLGQNnbNkRVj8O0pD3vrYDnq5f0YaXy3/8NiPLYxazM3rXeX8jelB8
3lJl4itt9zbfbBmd5rhtw82ZemHlw82TBQAjIXUNLHNxJ6vFuvnjB2m8nwM43QsW/S7bvj4uNsZ5
iFWrKNXRPQAuO4Q5inRpuA2qlFcjRFK/xqCGspRV07IlnXO7Mc+3sPnpwjcdBfuojl0ZAC6rusOv
HWLGpoQd3XX5pvSRq5KM+xoonA7EYUbjz7Esq35fZyEqbo62w0y1eB9pk58EUgceDdY+HLf6ZLtW
6yIzgTkMD+iKhO3Cq6LKQuPgYtOiZNm+PEgMeojBACjRby3aRF3GGyAYVDrdYBjBHB+PvRTWO1EI
yh7L5NzFoDMh4yw3p1nbqrQE9Twm7pLFQ5C3H//c6ph9abPprognlnxf8ibZ6UEJCE2AFJGjoKbF
am1nPlUsaSmZaB7NBQJpRguFUtYtEQPBn0rZXNj/f3u9yXHmZy8Gj7dZIc9zwNYNnUT4plCDq7Qy
LAI2d4aUrn6BmFjsLRi3gJI0h/Pq1DYuW699rzzvVvJF7V7d2FGZDb8DnTai2AJEzN0laOPpF+tu
9QbRC7bR33Dj7pSxbPdMd/avOiCCPxiiYcJUQfjCG3Bw5bzZBiW7qOvojERTescyRO2wPN48RJH1
45FrvDEmisQDiWM9Qbbol1jGeXpWugRaqYqBGKMJzRE2PipbefsH0543xFM8J4ayyB9yZtYKPxGO
RafSjWwk8bXMpT7onhuqSj/F3kH30zQV58YtgbRoh506D0taHJp5pNP8n2e1NHMjtODsDJ7gSzDR
kGrY1MIDSgW9nayvl4BsA5VtdgERCyIbs2iYvM2jAFpvLW3PKRulj5KlW/VWJ6YE7B9mjzs68jXP
GpZyCrwvNLQXs6wk0/naUDDtIslYqb6TqdpXBlRqiNTQAAZd63l69bRNcVDoZNJUwGowP3y6j516
xslAxaIx/O+L3YAh9YV7FTefDOsEcxYvloU+0MnNQbGJ6fJGuk/V6RXxAgtEmrAsxXvxWcc900Jd
viQDC0kkPJm+GtSyuRmc6Pg+9/OkVmYEX9kEp2pRA7rz6g+V6i8gGrTCMmiOd4taHZOYHhgrPdJ0
/tt5mYbCtHCRkkhuZVA+VRVD4XLKPouwjqZP5By65NlVQYJ6xHCZqRbmdtJnb53pbexlydhm3Aik
8qELrdLoo2qwjeJ1aKpKPk7YXjoGFFBWc4UKw4QxeQDthm9RRLA8duJxRRc4Vd0Cj3tr2vj+I10g
SwJQOthFNarbra+fLUuLLud4Ocdgo6ZgDuYezjdl/6HkB8lb1VYbhWod2Uly3MlT7ug3AskK6bgb
+ewUnrwfpVxN1Q42tI9jWMxuyUIFg3Fxmr1q7a5YhDMks1Ao4pw44OucoilK1lzkeIvsMqrWBO9o
3nCZZ4j7QFUnmoUw16kwPg+iZwYYvqT4Y//WNq8X8vi0N16avrlQ5CFMrtXYvpgX9tlu04x/zYzV
35QPrM9PdLOOdjrvS4YZHRnjU6+bDuVUO9m9uHiWV0X8AGc6JjBABphaZLwm6OKlRYAex9CCkRpx
v99/gzCPbXPOKvXd98PO3X62W6KmU0l5suPr9h9RDsum+xGCyut4ojKSBC4MdXNRHz4aEGws/jdQ
PmmwcPFSDIMr1CB25+/lOf19TUhVCyjSut8CWUqCamoVdxx8zwzvpVWLvOeX4eDo4OV2NnL9Rbfn
AYx7xyQW7d4h1VdC61rghoq0rVU9dX2cmhiEciORDuV4ZrFESCu5Jz8DFRWeewwOjm8c6XrdMMI1
O8TfD7PEZRRO9xAZX9igoebmghw8q3e62Zu1uHqDkLNr6TRwbPBjIyN/NtJuoGmhVjfEdynr554O
8hT3UfGWrcJ6AN3QLwSD+20RwJNisPj95Z4BS+HmABViT4CXPYStqhqUXD7hfTgwnRVaQTUNKjOX
3iPoeZD+2rdVdzsiBq67GLy9DeWhKe/yHeyDvqkQ1vnodeiajBkr4/8x3B5HHtsWrGuyGlj8jQxd
eVSxJhfeWxPD94zBXStPiykYLJcq3QZa4PBPz65mjTghe6wuQ0RAxPbYPl0eZON8fINB4oMu/h8M
9CXWHnD+2q7Pn3BcZHQRZG42sDErVVL440LVwb8KTUm6bClM7fSFUBXRckHyY8MOx6+JudwwPsAm
v/8oPERBfiZkEhURvnpW1/2298PIWKkPyB19Mi84wbvHv1CM7srRZ6JbsPzA1+/E3mQxZBk65X46
HNox/Mm4asxJJvdCbfn6scOklNkcciN5weT9so5m5MYD88HtpB+epgD0R9VP/7WLKdn7m2N6w9Sd
puRCCMf3hsqSkccWpPgPTPJh3lJx2/9dWkV2VqdbxXCcOWpYfICmcWubzMw2IxfWSHehwzap61t6
hrH18jqNfAlSeSdhKpMAK/gyS6QCEF3yXkW2WEOy9mogBbMXeHmad8OHrPzVhVhdUYd+OMcc9wXx
xgez1K6sNyEnui7UGVNBGcm3DHWo2dh6dyaraAsCaxhhlBz3kMisTLNGF5LtfRikfpI48yPi3zK3
PtMxNX3e5C+/t7Vh4H5+b+/B3Pi25P95rJZQMKXcPMQCx6RGBhtanDwVsSR3SzMz8GuufyPyTC49
/znytEubCMEzaC8kla30R0fTJIgUEy16r8cPanJl3pDILu6Ds21HlCP2dUQ5zmwO/ewsRsoKYRg6
TjjuAVKUVzMJDF1cVboPEKa8+/Eg0z9dCLG0tzXSHYHwrY8HT/TDMpse6pThGcoNKoQ68HiEXKJ4
BYut4BgUdRmGwC2cqWBHyID4MA5QK9i/Ve/sb5K06LtZrDwixxiJcgVQRcShWA5IuOHe+BV1pOBb
KqhWbPtubuB0Eb6vkAnCgnaCw98uQco0rqMAWpetXLF4F/omhFL8GEHqvPh0UHpBPmpcqfA94UQb
+AklrsiPt9BUiXAdfKbylTuhMzOh9uWrPPWhRupUAWE6Ha6pPZAE86XMX7+LFQUSd4s9VmIn2mKa
YKg/z1Jgr791Ew3623djuY96QZokcCXmJQ6ka3sQ+jjRn8akqDjEJOAToIIPjb3nsUQh8hLv5qSC
A+G37NRpZ7Wao40KbYZOAGSGfxvPhuv9ZGt67Pr6UfO+6w0zh8hxKQrVK5lYFtpHZaQJWh1KSUGc
mr8+pGQqPjoXX2c+wJp2TgUP0gt9z8lbhhhHLm2hCm/zbYXIftwpVDPb7+buitCD0YP+FueZAbhx
FMQHyYzcLVdR0pb60xR2dvM2TDELJiv65rkFylwW0ZKNq6gROyuIAevt+yAA67fVYsuUWzPNmJY4
4If9mlpMwqwkKcJKdFDf+mbS6UYCd2/eMaPI9knNcyLPOju5NOcAI9tDQJQ3UppdmNFmhKKBW/1v
tiCi8A3l0spR6qwf+/Uc7zmY2cZkbwQQwQeieraHBukMJ35Qw8m0oS0W99mp6AFNOnyfjMeoGcd9
V/H1uhFLfOpogmulD7i0Uih+e+F+zmmIQgO4wxKWCT7Fc1NKOtggGBdfK3WPNZrsP0+C4S1i6coX
E6Er4GVq6RS7NdedWRR6+TIGZMreA8AmbaiNtQMRohwT5NCfvxH62sjnRZiWFyWzMbFBldrjtxNh
+yCdh8uCX3nDJHRGN5foRsJVHWM1BKgpoaX23d0gLvGjbTRDMzbIWEUqypNw+QVljApK3Acus19Q
m4YK2fI/V8aC4MabHyODBSDnlF3cow6ZA1lGhmGeTMDTiug/Ip9buGXkB7coZrQmNaJd0vCzr5g/
OhT93CtjzAQGcYrOI4am5bvK9h/ee+kgqGZkwma7QezSL1V1oqFJPG3OT+3rTugzv6dekZS6MZDM
FKk7/Sk7XoHcYu0Yjaa/G6iag1huiIW9dYv69+Jcj/6NmmWm/gVz7B9WBk8qex63gi5tvNMPRec1
eXTtFNEnbwmFPi1jtQ3jK1611Ly42tNIfkY1XuCXMWEWi3hBQZgnAyFKFobsmPXFJDgIqUm1B3bv
ABMN6DaFxOXlr0oUXlUKGhBFY1Tlwi+JYbVdXl16n4OpPISUqpojTPn7IDqgvg3OKb0qs/67Ijac
rmYDuByloFwldTQqFYOK5UqB/weK7Bo/NBF5xCKaKdjq/ZV7A9Z2KhcescGD9MNF/1ZLB8K7fy34
oW48DFrfwwSVZ/RjuHHLmg7swYPcdkpJPx+xYoO2NsYoJro9WJSuRouzc5gR32kRIeUGL2sfqa1p
Pc3Vw/HKxxLzfX6bXUJ6aU3iZXRMJelPjsso+C7qgImSzRXxtuV4ASpyB03E0LkGuhyUqb4V5tif
DZNtfXjqSMEIQwGticiaHeEFL/c1SZLaW/bwVpbrtW0hMMj/lp313QTZiuExqXqCHpIHLcqFLR6Z
A+aybvAfa8yyE3tgZurjBOI9kmRQcvDurP4dpeGo1cClOlti9y/sWXJ58cLNjfHonuvWEYLYtwoA
srBhki3r2n1N6A2t6KgpXg0M719k3Y5SCSeCYmfqP/d4xU7XDdB+7WijBIMOgR+L7CeZSopjLe55
bsO2bQnTiRyrXz54i4l4G+3TydMXOfZilUsIvJfWsFFi5U1RRdS9Mz1iS0HqHo+u+gT5KyEIfEAK
cftgxvfU7C5mRZUnrSE8k/Z6vrm9LO88g5kIganzWuaTv131HiW7TEOvDgMD/PjQlbkOEO65uXdE
FuvFqUOZyWWFg6qSuiRqybypyvHwxpH4JbxNTVD34Wq8dulHPWv5LtCo0fSmpibPMt2ZRPfBXVO6
Y0zwgDIbqUiY7TVgOoi/0z1ETxJakVBRbWNMHgapmHonE4jSNqyZV5pw4SIYR7nJpf6OFmTNHJ8k
X1rwTHvqnvfcQgMqFajt5w7MUHhiJ2JMtW21xWVmTH2myRnWnNCtk+CnpC4SXDTv8HrBH45InX1W
wnj5B12613Or4/ZGYr8StW5TUeUS6W9lzuVrbNqhD8LbXP2DW1GBX3ymQNWz4iUXACmxH1KmnjiY
8UJ+kmskr5xX9EsD1rXiGQXT3VLS/l2D4tSuU3CYbJNLbY1WIxiHwtMZFCUBU5J71AFAyv/SXQO0
8M09zgiyMy7nTGqxGMO/0GsHX2D4E8M9q7JbhPIK+YtJHnqjDtx1CUQFsqecLX42qaMdb+ghF+kz
R3i5ueSTxxtoPUfnfmIMt+nQ6QzFYakFZ8qzeAwBoJf9636VAJwAXrgzj9w14T3LxywkVWSdZ59R
MsC0A+az4/s0SNm/k+uU8cBEN205rPQ6UlapGzoyhuJ3ayBuj8ZtDMNrnstzxKFyYAE+OXSErtUJ
p9r0okjySO6h1xVRWCo5Wtj7+9KxIad+JvUDQGM76xTdK+DTVvFDJ4FRyIj9yQwoekjZwu0jvBA0
SCJQChhev65BDlq+ERAm0WFPHow/Z3P/uhBZr8UI8F1nqxnrXL7pKhzqtUsoxC5hGlOfHMOqGpxM
WYOgBPAjSQvciqR9flATZRABJ/iRxn4GnCUe7UCqlE4wBa9bv+gQCQU9g9KM6wCDugb1iQmGSOGu
sQd3e3Lx/EZOFVDUH6dEiK3dGX2N4MyVacoR5Cjg/GODW4jpfD5guKezoZ46wg5NlhEZCnZGQPZK
yYDKLU4gLVbFs0l6+0lsW3TZ69BkUcNAAe1fWhcN8rXAR9k49TcI4Mnu4SZLYI4UIyPNPTDGBCpU
bRuhokM5wCKbpACzqcKSPiW5RUmnS1sdH3OjlwSGZfYoYJxjIVBLgfpz8r1+x2CO35k5hqLjUsi2
jg6iEePCPba56efzrNnHb704qotOgXY4uX5yiDquDNrRsNMBmgK4gHjqPb5vjC73M7onVHmqJel9
PmGuhkRCRpEzKXZn+iWR0TNcelA6Wf3URVdBhEExxpbZmoE8b6WAzAMdODjLba7hAiqLXCgdcRbR
UAxZBYzcmXHYruWieJ+qHx4ODDpVKKjxqtZvwTbQBkAeCT6N5qR6ZRPhol0n49pbFTjsJOB/QGrb
m8fFcwhGb9FVM5IpwKRPwOXLtKO/XPZL5C1DPtUaATMGtwZXc8u5BgxLCAbr0V5QQcKvNiVVR59o
DvvsOKFpOkwmvMCWblFMIFZDg2z//NSGfKHgfab/4gRfwyd1PgcZhwkCpYt9+lFRlGpcdWWi2J/Q
y42MVdfCf8q8V41RF4gPzsZVLcPNHPmTn8GvRxzLw1ultqHXf8D3IDZmIzGzOXyptJ+sTNciF2y1
085t+R4eNRoD1WZIgVd/mV7zO0zCJ8hfnZIC7IqRfZIY+Sf3HhHB9MSkX8dBvg4m5J0M2YqMeEXk
nOBxbbav2YjwYKM0CFEjPIJhMaE0kUvFh55mtIvAS+PN/sMdUa6l0Kg3RkFKQ7PCBxfFc0USmbk/
tgl59IikaMTre3oOAQfFokg69m89sOVQSDwKEj9UFGP7daJ8FPfyU7b92k9f9VTAvzL8HR3d8X39
Yv94BklXAsylq7E2sahLLw8KFP+PsiOvXw0H50nZlcJW6u0E/wJ6R7vvFmiv4iAAAwwekHQ4x7Kq
LGJGhg6ORICptZa5xw+2TI3Q+/UtJMF8sNDl1JxysgtXGqn/QBoZ4n8o1U2laPZSaQxQJbygUgb5
3yD0FJfmS7G/naVwkrIOedctNK1+D3ixm4fj1wlj5vAVfChev5f8UwOqe/ogxKQuUDy88YZjQjBG
aDlhPIJU0xpU/Qd6C1//oVP3kaq6nWiIpNPiSagLSDz9ry0APN75kLQiFXfYZa3Oiz2kILhlOoil
lnREYHUJINWZhlU0ag+/Q9ZVEL5JX4jQI3zWg8kOMPqxSMmLUMhdXRjXeXe64ulih3yshnbL0Ybn
XJUIXuzWa53/ZiAQR1L6DqmuvB2z1bLSBpf59JNoyaUkdT+ecu6fH3q0PTQ7MF8l/hhMrUSR5e8e
FyY+ux6l88u/nUKDIiXGu32RPEwJpItj5wJ/CUpcvyF2zkILkNUJSjDeNJCpq8mIoVbzEe2gyEv1
+PGAWv7jQrgyXXcYnJ/Vtu+p+81dFrvArQxmzRUJUsHCfzWjSFAjK8v0z6iB6ol2DIeY3Ecj3QGm
ApR39UE8KV4BEQJltIKf53od4+tCm4eSVCrKu/7WJncNJD6JH/lKats7ajhukMFr1p2psWAmCMA1
uAuRixnC0IGtujCERP0ZW3toiICdL8OZKP/d6qY7QZXvDQn2rhKVmnuXS1HYwMkeGRdfOo2l3N55
J2hpqK1774WMEEzt9gXEGt4IqBbsM/hfTP8peCndwAqEadFEjvubZJrbMHV3XyEvgGjHbug5K1GD
rDGqew4KSNUAz280T3HGr8TAZsVE4XQIiBxW5KusgdiB7SfDhBC0pfq+oDzhtqc3JFcfAcNlFqOD
Rdl79BGcvN4YDiyLIDwD92aXndU/L25sJYteWPfxuWJBWxTCwmE1UX5Zc9cVWMGM/j2mIbaZIfur
gefU4zZYygVOfeLn+DOdjdjaaTCInvNwIch5SbdTIISfkw7XxYosBYlKVaDBbnxAPRp3xNA3zU26
T0OM13jrXM0f7JZ0HUF0iAbi8abcm9aKYthT4jbv70FBPfRVhmgUb81W50pcJOpnTUDKGNYjR3G/
rsOhwbKqRT5X8KmiR0LQKkpv5P/L3q1VLpNle2an4uV9fi3klzLlEddFne8gPB770zaOzQR2s9h/
7+exzb5k8n4yIRNQZ0+z0Gdemyox5LaAIE9hYWGc1LbqV/OHn4Z3HihIfWHmSWRJZnHBl53V2NZ+
eBbUlTZO/gSeTj1G6oOhYyyQIdJSA/L58/6rhDNlKtl6R+I0Z2LKhOBIkjqIIp/uAUv2ACP6QxqV
/2jhh71+l0EB1HKQGCHAJXeFnOzYNFvsgildZ16RduCU97zkBmxjDfoO92U69VAoKXA9QnZG/ec8
cIPtaFEC/5xpKtLEmnfJHh1F+Auvefn9uOoRQedqU2ayQSwQzpXNQOWHSx11lOTWonx1x3cm1UjM
aGs2Z5yKHyiztkg3L2AT+iTjViorZQ3YZMx+WQudtU4QNxSptomCBNwqA0lueisbcwuD9tJS6VLU
iEtzJO8mW3BHMFVNoYQkn4z1HzHB0zyc76wxWUZ6XPMx2hi8huSAmrcZ6wmrLv3PT9vqtdhcF0qB
JV9J7kGEAvU7KCAKaDmXUk0OwMLIbh8BH3Y/fsnUXR6JANfIgO54CL/jc0bwLdZVTTIPa3xcRCiI
UF+WbLS0V8MK+ujZd+n2FcepLwpdo9YKBSwGBvM6kpnnDX9r/cSXOH42vWSQ+GsbI7AATuVV6iWB
J/CoZ2k/AxTBH+0k+EBQhSGC00soHNAMOsqH/bBe42LJCmXQkFuG6IcoMglVgzN7aWHVVS9kQO6n
YmttGXdN3/vpq3sNYyOVkdJIL6Gpqt+tCzmQBhX/zQl2skb5e1Wsv3mSo/Gs31+Q1SllN5/Tizh0
jlY/y2kB8UD1QC631OKTw9tJXOgJVvOV3ghRQXe/vylehunSfYgoiuHoRKwgf+msE3aqJ9WhT7+X
0Iv/cPzCbHDUMNA4TwqJFDqhv2Y0kky6kGTni4uPdjRB6CHmlmHZTxGAUAfKS4EPeikes3sKnXhy
l6Nfa1GOy03nCOqkiQ4BPLWB5QEJyzSwwPT52mu0FHUjNujcN6SBN3Hj+VsxfFIwCgKJWF1A0G1B
6r4VFpUQ9bakdw9FV03uuNPja1C5194hRQn0DWQ3gC01xr75BHkR9RcX2+kXDIcbbXN0zY1OAQWR
oxjmav2vfhI04VSPPR/nwrD/psgvNm76ly1qpyrKby4gGyOXTJ81pB+NGR2CwQO6Ar58SU1UCtTw
lI2Mof8LeBz74cp/96MCArl/1MQ5LhLBvWQs4kmNFPbtgBURFko8i+HoYBu7kucvIysYw/ywD8OJ
ESiLcO9FgXDEVx2dst+36IUS56Bfk0fyhi8d2q+y8FhF3Z7+0TRm6rPoEMEFTJgFegz5GeTU9iBO
lN+P3sWTKiEhqDYMRAQ9Ua09FYYQoYLcnyLAU30aoFGQlD0iihYu+61hmDskx+ovlAq9zW9sCDQg
sdbyZruZH0KCPfDigM4Nm0Fy1stj7zaXdaDPW3MHTcnXrZNn1sDEaxOUZ1oJivX2380wksTjEqSR
a5KLLW92JipYBrM6x7vdiWeoUgXJqMBaVV7YhN6iYwRMO/Drn5dR+pU+pfLhR0qODRJRFdUQbJ85
2A0AWhXR05hNM34ChIo/cZfYdUWbI+YQ9U03+y+YtdKigPWvT8/Du4dpNE+0M5cgOGT3BAjjwxCA
awlx90/k4rkLOJj68FP3XgwniEXaiusYXCAMAhg54nWMlLU17npnRTG873p3SYYoRwCX/gzoOLNg
TvUMF0ShpoAj5p4fdyevzmHuGYORGrRFy0RbpOdWpjibZ3nsChJOousZSzJoq0HaDmWIdTRbl4GO
lC58y9x1hZvg009SZC9x2y1CpX2exr+Pw6knT1dS7KiDqEqCI66MLa5JNzSEQy2LzkJb+w2D5U5h
UM7ABpPTpfyQAQC904tCMJzGznbY4Vz/oeth67DWSlVdiQa59EAb14Q91GNN8jHMjt3hVl0ISgnE
F+W79gdztBKIAc9JvqpELcZx/cRWXWQ3pOc+ikR4LwhOm35zPnLoYqOVHGISUiLTUw8xackkRbBx
e0QcUq/oO50gxjBqUbDe4QUciXwgp1isc6wA8fGj9iTmLo6Z3ZHbGH/qAnuCsLMY5vx8U7kJxbmR
lNQtCt3dP/mX8MVoOzQ4oWx7yRSkUVqXYJ7sjZ7nR1lYVAhxsLX4Rx86eATTZSc8GBqzf7vAAnT1
A/3sD6Zio2/QG3l5bGeDjunyeU8mGhrT/ID0LMCJ06FqLwnnPfbysPeopmyL/qovEC9rW0Uz9+YB
taAjtWiEBK/jIOSh7T5TRxh7C56SIIy+ZfnhN9QLTNroCmBR2qlysuVmwBi8sRqOBcjfAt+0UpgF
xL9rnUdLDFlKgDvXxQOA0tOrWl3CMjpZsSjg3rKZf0x40p7R3YTFxDf9zB4e92mEJ9Zgy4VUwo60
PF5Ie+N75AULVu5CAFfwmwYq1S0nCmxOoJVG+/tiHZuA/f8qCVtQ8b82UkcHyTRSD3GYv8cpLeyW
ghQ7k+c8E9X3rzLt1shmMCboB0x8FaU7gDsGKn9NRu293RLr20CY1Qz6tGvNbbeEyx04dfjuY1PE
DXHFKpFRkusx+cX8KtHhP7zAFbQvti5S2HXw6U93ku/d1A/PN0RZOshScPOt9THgGD4ydgsOhoCS
JLn381K29lJsZOPWre4e3KVtQ74vyTP2aKO0Hp9BwH3s2lSH4wsGWSZGapLpFRjzLaWluPqA8b/t
bKbO1HEMd+X/qJPRgn7tCoiwKVvWn80kM6k4Z/z0n1tgifUIpftsg1ID1rDpJceKIalQ3KggWdgi
v2QVmQv+0iUk7B2h5rlXTrAz65p20cQXF0vm6D+D8c04Xv0kdsHua2USc7/5S8O7JCncMyOj5rsB
diix3kZNqCDYBBf3hk3ddjAMoWyaqZOBS+o5AQkEgR61mtCx5tfkiQwRFQhsEBc3dlbVF33cXJnH
26nyLVTdAsQGCmBU4D1AHBXcqlojQPpl+TvhiLrEtxSbpZvqwwxNYV0pLUy6kbutRW/nTLUcuf3m
x4AjbUN4EmmQ1VIJkb+Hs1T12CZBdODeJXxgLuRjyPjy1XPXR60oV1aJGxqHGHSR6mkMVno2K9Rw
fcHjMGfUYsL/D9DfKxrNBr4q8AGa3CqNCIkLC+jE0+np/NkSeNB76tBXXrMDZbXqeG+BMcQRpQyi
Xn9XCPK1aVpjJVAoAhoMxBx1EzQLLwh4dcidrDPgWBRfYuDVY7AQPTO1yt9TMOBZIvNC4sktyXRK
nN3t5wanlI/781FbQeixnsY4jUqTUN7rk1Dg0SNDa0cJqZc5CcZ/vCGpplNPZq82oAfrjgtPaUXJ
/7HcwJu1I6CNnvV0/8YGdlbzbVXrZ7FnPskF3AMaJMH0ovCOUfcbeogeoATEAKd1YtdiV2Di7ptE
CY0VUpXNNVDNCLVaib3V8GIVkTsgmCzZMInNvd2q+s1YVF9H+YJhXxzQeQ0f8WjDjE6m36CPftZ7
XJwxiRWxUTOrzoWNyc6r1WBvVEuv6gHCOgYVbMmrJ3K3Pe+fDRwPBUKm2TaM1Ahxc7Q4BcExOiW5
JC9ZiVBSAOztY8jliINRp7jT1G49uEbM7pgYGHoRO44EgftDA1CdfrFos/CT9Yo/h5OW8KQ+PBve
gpVY1hghYb7lndVqUkSIa2IZb84xCI94ED/9z0+EO4l4WMBXmFOBGWmW2hWjI3Gb/+JnJ7+yqgKC
SjO2dHQq+MSTcMulz7IxE0eJaYXVbTU31fXj07Hs8jv/XbE73rw022Zz/G8sfvLLAWgVeVmA/6PE
X6N6Rv4B1XXDmXvwrLIgtCsTUvCRr8bb1LKURdniVEtooOz6VyQVs3zAQ1YNqdTyHCkk8BkhM4LD
OuNRb2bu3SE3tLyXR4w6gz9SJ/vnu7ALCkSPk2D0+ipnImju47Nm5Uoqc7m3SIXeIb07cg+H3drQ
Tbjrdr6/I9nRQXJ/+Zh5daT38BG03S2aBugZECap/bQaUtY1LQGzGIUa4k2C8L0AXtL4bzFQinwU
ZsbPdpfqYnr8EnUGgtqLtdpYX1n6b5lGPMncHMoUsUM2jDrJ8dhZ78z8T1b/CtrB34C1ZT+89Y9L
E/SHvhA10L//muIxAGP86tZpFl36wnBw4QVU64NO0knrqhtGfcPp5RsiKd8OAv/59pqZkEA28Nx3
vRkDyREbFo+D6h9Q0/qlF6uiXRq94ADwO+gZxfw0CqZKtpJmFj13Ly2QjLoXLQoMvWXLn10Gvdot
2hRhvdJ3R1tmsVURcqssFnhbV2YZlVHKkwJ3nkpqJ8ZmJAw/rIujKyt07Pg/fZ6ASjFBY1sXy6jW
0ec9LZC3lvpNJ3wUJgl/G+wOwKhnr2SCyJxUE7/Qb7Lzatk6VN3U2TeMQiElr/rXNxS7t+oZudHY
IQp4A46urlFNNOthdmreoAiY4iLbIp1ta6UfYGTOisntH2r/91ETPxZbI4OyOvzkjju84lQ6Lksv
K3c/zB0tcZDtVdYh64K2K1e/mxMutuFJ76uWLkfU2nDwxAHtDUyoqcnVD+3bMKbrv471YjRuD3Y5
80Q+8bUzCq7RyUiEOLPb6Sn8SXx0IJPXmxvPSnqk8HmaoTb3xIo/ESr/2Qz/hMZBSM0TBLaQCAYL
vb6sDFKWSOZVJfbUitnFsX9laYEhQfzv6+9ngYxRUCRAbdDaAq5kQPbwDkZRlXKbuR084Ie2ZBV8
PEHRuM2/1Z7L1CkTDBjtqkrsJ4FHuva+vLxzzibmaSXbhFNsHPz+UnxAa2RWTSEIRNBh/dGHJOS4
CiT1cnp2HGtZ6vSKh+OKqFS95G3Mc8KHZwRwusB9BwjMk19JfGiz5v0irupSjgvROZqm/jLbPmXJ
Fe3oGNSBvX4QyOqqgIbOCn50vhN+ttFUjZss/A7ERM2ZB//kEsDr7ekBTFxvgRyT8dOg/M5OTWZr
qOdVcsGcW4AW2sBF6enR2hPQJwKqY11qiHHS7R3MZuMUQp1rRfOZyT2sNzg/hS5vDu3dJqMD84XG
iS8b+nvkS4rPeWd89U53S96uWctSuiGnIUSsfYyD5TWWW3AaHTR2z2B7HFOjCTh6RXXHMCCoSbXZ
LVICemPVPnJgQ7xNNSShvFbueOKwZZp3gEyMvJhGOR0xFrMUV8HOKsY1KMGO6q6d/yVPx+nK6Gz7
bjDxw0Jog3U2oDCVFOqRACfPBLgvdQzYd+vU/ItoQQH/H5x6IiNE5kOGeM/EB9IPm2FqdOfZc0t9
cMa6PVfsjH0Zyoo7mn0J8EF9KACmSwSQEKaV6oqYv3tGGLwpuohgF3IHfCoRt2tFz4rnWN651Z0Q
Z8W1QSYTE2qEEKnyu1aSWNofteebY0uZDC3gTJ6fN4dgsW5AhHnFcXk9jLdtiiVjgcESdTfbeSMF
njsHODhjgsE16u01277PfVTHlBzV8QIyLgEOkCJY/m511ztkF7127sqSrRIBHZbdxwMbH8/10OSH
6ih7VW5hEZzEZ4RdtSc/sBkMn8aBc2OuPQhXKC4bn77RGiamrPYqDBtcrS18H6fVewY30w39jBbb
8nsZ6hu2T3EWPfCZRddKy0VabQC2gWrq7OzjNDB4+Y+cjNnJMJp3jRRtQQUW11MhZ6YntB0k6ZFl
HD9AOzpo3Twz/eUqHMJCNhQKZ+9I5yehiYN36TmuwHNHJldKfJJLaB/l1uHHyhfTEhQDR5ntgQps
Qzbr8xScwrM63Scr46cx0qErooJJNDYFKVbbRzBucMg8d6iSKdHXVGEvvkN2WyQcKgIY2eNEtq10
9nsd7CwStsfg2wkPFZQs+okXPsebBGLxac82Vi7g5efUIA9CtPxbvAzLq0SaFF0vmK6mS94cveEk
RYcVFSzd7rYmanhDWFavqefOmRzw5oEUJ7Z9BS3+MLQCTUOBT8fM2awk2BGamN9igsrkmo1TLMGO
V78uoMFs/K/AW8Mi+LjCJdRxr1dpo1KlQuRHi5eqV7cyDWcv9f+ncmORN6Ib/rne3i2ZZEPRKGjN
OPqMOzlEHxer8bkqeIW9Tmq0A4mzNqAFD+vP3eMDL9pkS9jndth1cINq2xE1RZr9hsCTM3Xcu/dk
xckhUWQXowlb+ta4dYYSMWiRgSuhsuWcviduHEtzpdGm8GP7ZSSmH+ElzVG5bSdyzO8kcoEPG8ha
1/uEayPghMVXxoQXcOFKsDk5xqYM31Xa6rcxP2hUoVOfY5zl7/4IIGALnVz8eBH6RtLw7kRoXS4O
CpGIKpgmvgvqJVNuNgifxFBwQ6YGAxiJkMtHx8WgqJB4dFbowoSlZ31iht7E4DQvV68jG67zlKKR
lmp+TXjhJ9BGJx7VLQEQMYjNJJgqHZUk4zLjMEr0G2iaGSmOOXJ9nNl6UBDMAOmwObnahSgqvigR
UN7J41WNtTcv+xFuyuJIqv5dDJx5ht/hcFL9MT/357FtP+pBX46FvrrVE8bE7ymBaHRWfnb/43Ej
EdQ0nWC7Hm3SVPmpoG/ycuBH/+ondtYbuBROYMikXqtJ4YayG1nW1gLeVoug/8di8cCcFUBZJ5iY
AeV/v6UMOYAb2kauKsZlA2PJAer03dKpvQdaYcMjsOUPVwLuFlZo6HDKC073ha4S8XxMYpzPrEe8
Qsjr1O/XgmS8rqkMgdeL2fburUZM+saWVgeeumpBjHgyFP1PsaUPoV2OWJE/jaJXawzpErFfSgub
WOSJssExE+W5j9J5Dr79L4vNJN0jHGtorAPbt+GceRHEUDWevW/3AGbVNG0qt7vyLzz+1+IMlxco
DmZchHLttmlj7ZjMGkl9vuFnAYyKxlMzuZBfwV68eU0Xkgm93jNZ2CItRPFnGqrfNq7PHvPQ7DQ9
4liYxYAij1uXVLra9qsqVd3xXTzCbUnTdfvSUiSHvnPZbIPqpeg5oU7KqStVqqoPtV9lOp5N/CDG
1aFdiofok9xPjPfo9DB4Hsw+2qZXIMEajyJa37iEwqQDCtE2XQ7tpO7NkNHD2XJfCR/a7aWdCLyR
i6XmnUqk3ui2xJBejczu9Yn92w3E5tiIHFqfb4b+KxluscHWuGohZR5rNVU54plYWBM0KCmf2XF2
brWeubF5JIOUD/DXls+6tYKtLSWtugzCe9TZIxc1BnaSCL2bVTChGfEWHRWO3laswUDV4D8j4s98
A21OqiG+kG4G1xsG3wj1Iy1eDUWRSM11DE3PufNh4eN05HNZkHNU3JsljzCQVLiGgOTPCOn+rx4r
JA7fCLFHMthTtH4VPiInvVvJJKCRLbJ+L8Rgsw25Fu2TguDTplcQ+A7dfll9SGRdeeb2lVGJR6Mh
NbIksHoEcB4kCn9VAxp0oqC4NEU6cRjN86/hbyOrf9kzwoso/Ae5e9FOcFPfaWtN9U401tqgMuMb
w7VKZXimLtMl9k5tj0wZGRgapTsiJ/wzFjLgLRw9NsA9L5GYGGDOVKwjpW49qtJPKsVZj6LKFUq1
zH08hhRS3lQrjWMsRPODEJvj+o5QSJCmVSaWocwbuDBOhgqopJqZOgdnAJGwJJ+SKqG2wxVBuS8k
pv8Vd9qqaPA6yyEmD2LJ0QZe6fpJfSg3lO8c9NRWjHHcrsgtgl87vcdV7FUQ3/QsE6/8oV3QkGVL
c0G8VEz84pFVZ3j/G/2rxNEuukM4DV1IEAfyZiypu+KmCRZqOKVv+QEMnXSkiVqmzsEI8ujFVN1z
+v+3HQmLV35Wt+lt9pRWfDOsMmWXWcThBHCQlXSveeoAgcNZE62iOPJiznzk2+X3YWqdmQkk9Jkz
KPxUhnYf0mw5KDTW07ILpT/rXLIiht9psNDFZVdH8hmPoSCi6MwwBVBIsGZzE6y5smHOjYr09TiC
+aKOGM8+pqyrx84+4vo1xSZ52dDFH4MtGo8j3TKqYusbAh3PgnWjbL3DOhZE/DSmz8+p5yF/rMPm
skaW2czR/1oKjt9sRDaBYGEY4D1nJkgOO94JObWQC8uu61nrJ9PP3Xhv4KZt7RDuSuXdyS3RAygm
Sf07FAkfvi4V49ZfYjQLM8kNOrhLWFwpWBrmo5UCJBDWIGxiQsCrfVcpNctk2uih8gS4wAkBXXql
+t74N9AfeIglw5veSYnBeDDN4mpFtznVosefD7kwbWj/7uPyyk5PUIGtu9eNmVWoyEb5bnfI7Zds
lEMFTLa5a9lsUiPSqMTaDDvEcX3hDKwEE6CDSXKPyNctrmmStyvvtABU/hpYm1N9ump7D6EG7iU8
ElcaZ+obnOUYY1hyJ91cD2eUCZzJwEfFHnEnht0zva6Ex0jnlTa8rK96rFHB4zuXBtRJ3n0EmJp4
0S2KtrC9r6X+24ybZQ1dA4yNPel12rmcRzhCF0diERzNv4jJooYdtTsfOthHlkBDHwxKv1owDMIQ
D9st41DepLzoe5p8SlB1q8cVRjOA0YwFyd/VyoWHi64A15k0dg+Th/Vo8/kkv/b2QUiLeh9fbE8m
sbcyAuNFQg7g+mZmwf8rWNCf24tfVtNo46q+W6XBMfHt+wFAr4LyAb80ZHT7nhXZHUkw3KAXlShW
wj5p87FF5+4up+vU/4XkT10nh2hjej5RezJMTjmMZFmFD/4j5KzbwjTToTHZmHE7Zh/eypdQcrEK
wxVKNyS0lgeJuHeF49RRN2LoB/an/bbAI+7HIxR1IOjqFWd7pomBeKPouEhf2gXgCSzRI2en0CQ5
RLGUVuWm9R4ks8gWK2rKxFx6lIDOpdLeSS6iNy4d8BEdnzfKOElInBsLqQSaY+3ZgtrYccVIrX6Q
/5wJJRRzWNAbR1mrgLOhisn3HPbR+UcTpkuPtcn4YF8JpJeTLJyHcbRyqaJ7MYyT201aUlpJfg+S
TqLf1Wte/PO3PDQJ6smEy4LKXMKurR2crHSkzdtEZBvea4E56wgF4vFkpGJad+0csn+FAi/C3aMq
FpJ9pVj+5ko0nhU07fxVsM49UT8E397ljxr+r8Z5AHgv0bfryHAadk0f2/Yk7wIYgYVeJjIZK60P
VfZL4z1Yrk1Y83Hy4WktY2WY66/ZCXd+st6F5VZuGJhJBtTf8aGHLK7mOikgdVoZ7GSP8QPe/hHk
svJqmK7xH74iG3Vq2NpTG0qxtGBAy5b2RB5vFD8TJqeCU702k/fmC8q32zWs4a3YqnTIwF5otS0D
6tqBJEpBNpy1Yrq0ZOd++jSn+QJpa/ZvU0btxjLhzwzaaMN0/hioJ8HPlmYWg3kQTq45WwB3JfE8
px+eNeb+CUjnpaDReAz3BTDKFnvbKZkQEjoVYMXCeskW44gggkPlM0Ynkpmlu37XVrRfKqOk0slV
jqbC0yBAOqrp1qGA3n3bRTUxwoIGOmG4IHhncZlr/48SMg+bz2YiKY/vA+JalrNg6ysvhYzoXC1u
tGOfd6SsamJWfFxjOnSiqwHDBAVoSOxNKhLwQoMWHqtHegUPTTdPhP+aEmz0yazhhyd8tLqD++KL
hRc/cUmteETQ4fZCfAQuAbwX+FvyXcs0HIf6Q31wFzX6fV9AACtTZCN5ms7Fu0ROTHvulpYKD+e6
uDJZ7fBY98J+HXzRcwrPAzgckrRqoOowOL4tWIfGSSLkgrnp5cbmJxQAog3aj3JINy/mIvDMe+Ko
RYvYx1Z6/a0MpI1Fb+eqo43EJA8hdxrlCYmiQ/OUrM0x8PCKy3lVoMXkt/iyzvki5ZsrVRC/1fkA
PmsOGlZjNwcNUSOEHdcyZsz+HfqPHnMgjiDYLoR7ggdw5+tjPPM90SlMFCF826xmrkTZehtxLW2F
BSBiZoTZ0VTdPwkBvBwnQGdCl0fMrlGz5P3J+WYvJMgzSGG9Ste6AWdip8i601C7XK+5fWpN5uQX
mQmXQ8Me11He9B84vjipk1JEICvY/AC2EjsX6960aKWUP/4GfsVbwLIbhIZJMHgvdEU4Ju6C/V6a
UO8L0KpILWdWFytenDHgycM2I13fzAOeAdryNIfbjd4wL1U2iAlZ+VLie57RSO71L9YETFH5t7CA
4v9DBaWVvZ7XUYNxjCkZQLEUFvRMZEz7GdQyOF/zzX/Z5d8v92+yt+pnLTS2Bs6rYNtiINZShBSf
mQv6mIfXnDjbCnxcO9nP8KeLOV/gbUWkDUi/hqNSWeJJ51nZ6Dhj80F7dYO8zjTok8Qi2PN2lo7C
x87azpW00Xi2fWqcRX6d3BGg7bn55Y98dsw75r0b272gbVkRr0uznG1jK/uebgtAnFr5RT8HFpYJ
CWRh2lRlUbr3uwL39YI8ahgYcQUo0pfdVz0rVX0k45FWWwI0RGPdxNIlwCjpTxduOeaTRE2pGNrE
MRFsmkQbv9c2Xt1564kYst4np4CynQsRMSqHxYjTeAyjOGngCCjoWLTAh24FgZwjJzPEqWgSmTwv
ZztUC4shNZ+87cCLYL7TIwzcHNn7xq1mipDR+6zRJOK0MW3aVaNgIJ3xIEf78fuhyb6IERV9Mrpj
r+KfO8HTcQHpXmGKtvrqKuLuxnJWA3HbYV2EtsehUT4hpkc2TcQSQSIxHA74q6lHgD5C4K66KmlS
/wwQC5MWcp1tZXHpv3mZ11G2qMRtsm7aXnaHC+UCg3XW1a73NowEbaXIyEcF1H3/Yq1SAA5g+8zU
XVX2vtXDVTZs3K5s/9KJMVvS4MzB2PVdh2OD4otkBjVgbu0xy5zEUPpmxj2HvxMN1Qj8rHGvhIUe
EyUGFfbbcp1kgHVN9wZ/5yxoZRyWs6EEUR6fzlGHKe79XHxnGZeQHd6RyRFwnLUkPi96lsLXbDJ7
rdJ9twjaBSHnb3T0kdlYyDx5fdgvy7FOt0MZOx1ufYgm2duuqQgwTrzWtmPPGkR7PeumZNdw875b
XSXATRmJhnafDxuU9h95iu+przbyLcZoyBR2uzBvEgXX0hkTKiUn8DV1/KPG93h2aUrffijdYaPY
yqQf1bG7qsyLuDjKKmAjbkFXuFTEFRvrXTwHQW9gGaopcv76Cpmt2mo6VPSDwTt2ISygn8Cyz7M9
VIvGQUNsHM97qtC6bDd1Qv0rKQRr3SD897/CgYYJvTJt5i9a4O3yrv3S4JyOn+rsW7g3Gsu6D4Uj
maRsPKyxKstZ0jNjLjIILXtlcJXSmHh9CXQaIHAEhIbjgyEig4YCZuEjA46wdZqEZ3CHQsTXMqDs
poZFwO3IUgtPtXR29qHpAMtNSNcVlV/2pkkfL40dPyLOFC2W1xY6JLR7BlRzw8tr8YbMEctTYA2P
pMiyHG9lVje+H8zGtJhFWBZRN+mgQN5oD59Kykj4CeJGJWTBTrXGPu0WVb+EWxOPbaN91LzHejxt
s9YTYUZy4L/ritWgazjzk30l7qPYb316Fjb1tbPmyxD88hqky0GJJLNdZI8itlUrajx8rrCsrfWA
80YZJKWWBKoh0l4rANiBGOdpAYEkvDKSMBNjKEUPG92wqCB2n4cuUYsPrmeXDGRFfEOqxO6+6Tgc
HrqveItgA8s2npv1lC+jR8/+CYqDnGibVsV7V0TOtHUM7pijsdxnK/SitqjvLJUuUnrSH5U6w1jO
l8h9/QVofzBQ1Fv7JtiP4P9bN9uE8wZXF3Xmjb60sGgy/wK9ZEGerg8HrwWNdOcRnmbrYn14tGn7
f4S+4ZRrNrRCsi0gWxE3hP6dwX2y4U0Z3hjeHrFap0xSYYEMViZJPa29Nli8XqQW/OmAnsxk2nev
7M2HV5l65AfBOy9gZZhTxRROEEX2DwCTun+TXueebUhfxnMfoQg7SJNuZBYxyRBXVroSOdMyF61m
yCrh0jKZlmOKsCprutq76AXS73+4B/Y5n4q+iINb6hDdU/XFqPy3G/vusKUKSpZw3bcjb4jcWNH7
5GwUrO/yNG1saFK56GHa7hFeM1OKdbbg4WluHQrLJ6RN9tvu5CozlNxtHT7T3WyYk4fyY+OEq4Xm
WtKaeSMMWhocX3NFtRLrVFTdtb6tiIK9rpWeG+tIqmoItJ3tFKC54UUDKMXkSNzOMJ5BiOzBNMSb
ysrCvCSneI/US6ow6bVf2wbPNt5hemMryNWyufisEFEppKz2eNkL7QLomMpobJRsROzROiuYN7RH
KNJo6XBlNC0GlDXR36lyonmcIw6ms9KSmP3j+0H1/MbUw5BPP6XLioNZh0JUYZdetrz9/N4ZZDl9
wFXvHuswg/SclznLgEIR6sgeFjVPKa4x3VFnH4s9AT/IEzbEqgKU30ElT3rZNeBLr4Uy5JOIYbfK
WpIB2hlL6zE4q5fHpkrX1InJjJukNPWKlWHm0MtLYbMT9Tge2kcP1p7a60nRC+1DhGjZW7qptcS+
kcBFj7PHP1IEPRzcRBy6iDalrS1561TyNcunQk7YbRhy2ArBj3vo8QnoDr34LrWYbtEBJrORc+sB
FCTNnU+efw7AFxWXgkl4stEX0gvFHWVmevp5oMKXQZIAIGXJdj+6i9+gDea33e1PlNMu/0JqdRlg
QM/KpH8lLlfEWP2PzmSyifdaaNROPUX07FZo1tvuWYhlcOBlWBWLI1lUcOenAGt0iqf3fHvZQd63
cUTynH+WNURO4LwBvAs8iTKvqbu+FPXLwrOqSrUlKsDZSjIe9SyPtHbW3eQpshctgQoGc63rbshZ
qXn95ZHZ6sKO4ilMzGgH7y+hq9csnLL9Jji3raO4pMUjCnyzFA62CjAxInCDaaDPNfwRO5T/PvsO
B/IZ1uUhuUUVyXOdciEaVNe3JZIEOmgbC5ab6dgOXuhrh/gqwqCG56+6Sb7DgsADF8bV6JUMloTF
echQYSGJnqu5qv09DDX2sD4u8AR8BQ3L3Pef9dsM1Vw0B7o9BmZaTFMT7oE8JqgNqCTFyO/vMZc3
ZHgzNHngByOTjFCkPeBUuP7vcMpS8kW6YX4KKliKxp9nK1eDe8LV+Z6RlUaoeluh+vB9Ua1Ipr5/
0R1QkWfbELa4UUjGgLEiI0Qn5DBUM1C0oxlximtE79K/1bphVpzlprZYa4F6blK6qqpDkoiGqsg6
rRfFKcB3VPw49W/76ddpLuNM8nvzokhUd0V17VRGcN6jHqnwCxAoiPtjbKXwxHvEqWy5dmlowQe6
38MjnNN8hw0AdzYe+PlCMEbMfPg0KOEgmE/6bo1f2u3O7fsxzI7iQYjTyWbY5tKMqmzctyo7tEvR
osq5HyzfDZf5D2JJLh0oAtmuFXE77jv6Ve3T47Du6Do42DBvwg651jnbrueFpA+6gOoM2DygFCjF
vYy5e/e1CLXbi6Cci5Y/YXokBQlZXW1MneS5NQJGIfxzDzo+m6nXKG95pugOrV0O6uaSarMa4GIU
oFBh7zc3ejgdW7g/gAXf8KNeKyywdcNH/kcaFOA1eISEBpxbqzm5vACQTVOvQVuAFoOtZFYmEIKv
01X5ESCr+GjgViVwzdOTMuCtCtZA55YsF4hsGbWArSohNAHfhpY9W903t+N87T3fhkyvouEKJSVE
GrkJO0pYet3Z4Cld7nfhaKV10Jxu7ke61PGdIWPjAjFpgdpXnCPtLmY2yJa5za0+n4lv0asXzz11
vw0F0mPSDcFnlqwSgheyWVeklLOmb05kA0Zk/kl9Cc8ipSDw4OE/atIpjsILDg4Fthrr3QylOTJo
0cGctZ8RyBFRCdaCpWjvQn0+IAbhB/qqfqW/gVj53DY5Kyz3ihZsJJwSba/VoTZXIK8BLa4yvDWv
al+qjd7vBrlPZXn1fdAMVUrCL0QDXAMMnbV29OGv2TGfZjdrvQG86gU5glO5C/lj1PgcwTDKzlyA
crWstLwq0LLdajwZT/m7XnpiXf3KRb/crB1U+UbUpeemWYzR8MMlByIKPhaWna8hHXtxmKheBLF3
jwymuIIcYkGw6Du2MrNXkLkmnTuF3Su3991MCB7RpQdMnDaw92jV8XQjYsxC068409xqqh+ZqfUH
MpfJQxVizbIOa/X/9K1RoPQlH3GK2W0mbhWN6T6mcaUfGGQPsGlFSh20RkXcdlm3UKUhZ4/UZ9Hk
pqKNR7Z0EnD4pkZR2DWbLlGBdrphiB8Tw3YVEN258FDuv1qAigl9u0RIy3e0f8wsnTct9Vrb2T5t
WTyvy/UEEi2c43fABg6iTsrwNSQFs/qqG7LdKFREvBoW4xCZBpOK5y2eh+s9z9HqFCYz0iFJ4IGF
H93KpAV70+dcUFdj/ThjIBTQQ2ZaeklPVjXz8AbRp2uIn8FT+No9HXSOu1zQN2xp7argNXczwL0X
dLbewDbvbitbg3iy/S4OWjns+tvm46/wLWoXtIaY0gAqPdNDnLctQcm42a8IaaNkoh6JGD61adwX
yYQddh/8jABut/zTlopZ8BS0sJTCDUwFzrGDbPGsLt8QiaIDwl1q2VTvybAOhO717/eCXUfRhtQ8
KdPE2/ZFPIgsMgKUBsrwAKQxE5VstMioiaTasM+cSZmXCEn4vyOqCHYoCJ8tTgzUEoZKkpLqTpLk
q8r7AU0+xE+9eQLh3VfizKFj4+GTwBupREN8Ow0dNRXzFOi/L7VznK7OQP93wQerhXG3mhipFR6H
hnUIDHTYSkamcczzCs4MMAqjXL7Irs8BazY7nlMkC7EydQmjYQ3JwBQ+8Abe9Iw+JDcqNU+dp9Jc
Rt6Bfz9fxH63j0wGOlwfxN7tll7KAiZwBdFAjwDX8rxpnoGiW3P1Bg7hlw7pEtQC8BmcMakUnO28
8aRcFh2AFY4Sb4dYxRIdOmhVH4KaAlEa6JdsJvgyAVjLdQz6rofLDKCXdh248HuGiIB7IvfvWiGg
r3Kyt7J9GyN/+blWptvsfPk73X/FLk2piLPCIuegySBXOxye2gsSkhlAKeMl8G73uuOIIXh92z24
yjVI2QRTHyaC2dwVjFq1yOQD+YjanX+C5Btkvxnt3kDak1n3pEPRBMjPWT8hHlJct0oU3KdtA3EL
10uDm1V2taDUetjr9R4nrSvm497KNgiMiEJfbvDc08bzJ0htLaZLHvMjB0dZkV08QHXmKbqazEOv
yh60tDmZCFhvIilb9qtD6KjbV5Tg1QsnzKxPrLjEXiubq31zE6MtJmD1FlJiwP0pbj2JAW5qikx/
dD8le98ARQO26TpoKi/QnwokhEHFiKq9k+6y2/LWlmoQOHgf6gvJ35x4tKLKb92vVuWJwADVxt8r
cbikeqsOfnIp6BlaYpIROcWrDAZ0iBDckuypPd7HBs/MHGgFmIZ7+HD8RCMKZB2jCg8FuWiUyELs
0IYvQ5PagEB9QlMfYkSNPbzlECHxizwlxaRYXwcasIVIngd1fCwvdyZOtdh9+cSz2+lmAChE5mTG
Jaj7Nus+it8MMWa7+85r1HAUREpWcZLgweusMyINEAn90ku9hKgSnk1ZoQ13pJmu44zuP55bbAO1
w3MZqndgwOmFVIdsmfomziaeZTYmrMC+6imiO4dVMc/edAfm3c1/6jREFjY/gxk7xMphnBwF3MSb
NpYFan8P2jBXz5i3Uh9eA5EgPMLlYhZxMdIb5BAgsmIgqMpeLU3J+wSs8ZYwyIkYF9Ocg3ov+gYC
ViwkPVS2ksuZ/867Mvpc98XbnlX3YUi9nqH9Lol7OpLzeU55lrXktqy8Bjo63L2+Jrw59CXAWbZW
pRuvb0IOA9U4wMxHQ4LsJ0v/0uvSVPH7Ghpj1Wt8u4KSeLWa5oabRFlWPpp+/Jn/Av7OBzYo1fH/
0TbrxYPSfVNE0Xz/bPWwxMtOSci+3Gs1rbmQXx2zqxIO9blodLYwFi9AvogEyY/32YvQm2jCTqdu
LJt7DMVPspQr2JeEYsyhNje512bE0uzGV1aBpiYDRX00Z6C8wJCGn9cKYUB8N6C/2PYaAE+G3tKu
JFBL/eLrN7SEo5Qi/4J98BXEaXHGit1d32/jau5mAdc8rGXh2NuIN0h/M0+Ah6vx3zc8XWjJZ/dD
+8vEM5WBb6pG1KTL1E1Iirv/1XqcK5VYtEK4TawKdiQ7Li0ES6Z5xSGsOpEKBIk+owaB4DBD4Wa0
BmQZ9S8W8Y9+swVwvdajm5fnO14T8ctjroN0B6K+XOJWpcVxjdgFpAIakEQBW7SX530Tvu5P0g/1
tc5cBJIEQ4aB7Z164kJG/q/jeqQBKri032HD9h+KbrwHROZ/zuvsC13UuV5LOXZdF6AZPusIpvnE
vOShkMqz+7ofsWlwmpAA+pBushTP2hpy8cafvZT9bQu05BQ3+UXYPs1ObORGL1lwIXf4izaDjZmU
97shC0hFMcbQK03uVYelzUeAzEcr7AvDd54Oic9ztmpJ5KMd0DFWXTo+PW4tjrn0HTOjQaXWkepU
5uGLYpL9DF6HTMijYlk28xDXrtmI6twIQuyviuIcbU7hDDuT3QzM+qNdrcDePQoEFvor1X2AoFBV
HgGVFuJh0UmdOiT2TWnJtDKpIm2u8hdagDJOI9Ul6dDvrQRuMyqN4kubCszGZow6MeX3hi+xsM3O
NPvizkUsS7V1oliixdma4dZ5t+oqP7Ydm0ZYRkzQsUuD98v6ooHh4DC5pIy7l2DTi9iT+Ic1nlCL
0IBdcC4SitQ6yVOn2b+Y1//QqV6ickWpoRBImnW5hZFcszejLehQq4RjcSv1RA8g23YYbXTmS1BZ
VOmZ8BthjAwE8Lt9gR6aYXvqcmQ+2NDZSTx1cJy38gNvC/jyjG2AQRN8NT+ezzvPNiZAIBoC/EqA
ICyzLYBBzDsz5Uqb+ThBRnvWnTQGmryGHb0sbasqQxwL5cAI7R2GeWjYX0+U/xlrKEl6nFa0b7Co
NwAA5V7IjYdl+3NY30VukJ1DZNqNcORv0XPAuqLRT9V3cnwvwb9xi5Rx0e+NQvztPM8PZOjVcZPP
ZYI1uSRua6dcsDCg7KGeePGAjW8j9gJIosbDB2WZaE2BIARM/OHzbkZgbM58mPOoRPrY9gyqrO9t
JFl9JL8ZzdDoVdoeCvzmuua2fPd/kHLdpycv3itHuXxlzKiLdgZ9S9gkqKFXxMywmssRm17HZPXJ
Gb3he6XM80M+Q0rW4fia1pgBD1sN4JBDCegptw3muPWk0Jp86Seg8CHnHJ8Aevx2F1tPN9HmrhUE
UyNzs7l+I4TtbYUXJV3Q0WH/styysQc7rtIciE0R0j4IjZOs3W/qlG8/Bms9BId+k7+X7SiBWdIB
UWjLJhEcDZrYIQjWH1/ZNwMJMMJHc1w+pWZrcegAr6hvvs4Ye4Md9VCzlmGgzywpXrgPDv+I8sIQ
wD/e4LUnykLwWhqF6IIbSl4zi5U459iUvoPavNGcEdVSA7GmEpGbbcLlslRv5htYNJr4Cf7alfcG
3i/mSrEPJoT2lZoB8fBBOky9ouJQ8kNJcSFbcQZF7T5B5OV+r/xDdtC8CR0TXhYQK+FWwSywo2/h
u20MqQ0OFpEVo6oivvAIE+4Hdrc5GSnYlRpTh3SQq+qkgiR1ZGc6GSDVPRz5LhhxIg7iv2cKMViB
o7zBXUVqbqi/4iIaxJvDvDrYJ2DVhc4MbSkb+f9ARcsLAD553N9U95zs0BKPKeRLmXcYaM9Byv4s
0eEtjK0Y4I6aMkj1VAleTCTONCMrCtZLTaVMN6it2stqYshrhIbM2wAAm+PSdpPj4IAh0W1JtiDA
Z7p/If6cn7rCS6G3L+Vy7pbHrVgeJ0c4hmElX/E49qrHlcM5WIpWBEnW3b8r/Jczd+Bv8Te+MYY8
0NWAE0TvexkU3QKmR0Y1A70G/ZhtIBG8ObrOQY75OgtsF/QVUgloKuhV+ASQGrwLBgFeJbJuzWyC
uiMjHL6Je4a19Ppj5p9zkHhobNLkg8tFMG2absx0rwzMy9eI9btEotwp1fms2UBhwkjKEprWdGR4
vYEs6hVc4/8UbR+GjG62e9DtsCL9Xt+AXG30RzhuTCLV4vqkPrVRFLS6dqAzB9wiQpDy9HH1ahGr
vYFWK7Rsh2N3V/nnOH9XkalvDYrZrFiAO4tgjENWjJX3822YgvyUFl2JF9KlmFPQrLNZMrs03Ocx
itW4NpNZjX211TBplGZ3btR58uqoAelRDVlmAKnwhQ4eEcsu37QxXZKWzChnv1ebhbyQNamPTtjW
sfjTgtyAEUXonwAjUv9CPaILMtd2+v7a2Rymy38A8OzXrr592jtp9JK+wR40/ewZCCmtvOZfbe5L
9LazPqxdCx6kFODKHMxE5JNqm29L7L154xPor0w8XfOyteEyUO733BLUFP/JqCxa2JVHDhVHEZh6
BF7Z2NDFwsEibj5pkytVpkDmml5HQvnbgeRzy/FkJvNMQH9jJJzG1yPXNC7Mu9SSkRjNGpDlYrEF
co8u8BWWxpPFmhsK4O8ctcdQjrib5hCh6mBJHGeAfRouG79TPQvPFzvDlZtS0mjd7CK2ZOK+OewB
MRe7QWWqVV2ifR2P040oGIh/QGkmzY9fC3DRCpsv+4LrhUN4Byu3Bp4BwMi34Cc54/W3hRB/3VW8
Tn7rtn20pL3rtVhiQ4/2Yzd8lzyc457p2d43ZPb1dgJAmuHSwVD8N463aVW4pJDUWgf/tmyZSR17
tSn89TyMzfy+ecfHUcAQxVl1T2TJBwcY6DDd7UhxKDkNBugX6i6ofPJWY86gMoeciZxCj+cgp/LR
fVE9lM3T0dZleJpr+AlymSWkpYHJGNIxZ+kerzRymlrpWXLViYV3y4l9Gu+5TiAr+oASIlxwEA9x
Pitd22DFX7iHndsi+5JAcWQK1QSmI8Oz4lU/5izgzBrAVr0VbL3+Ixqp5XxA4HHNuNgVbD1UwLev
V0q/ofDO350VsTtzoZmnfz+Y21TSvBtJuIjMhpqaVhFnLXXFb8KHWyfAUoL9xM5liBYz07Z8vstf
uChm3WCXPEjpHJD0S+bU1Zf/k0TPMfq2Sud7vhajNOButoQqU+y7aFZzfKZ0mVDWPIuZk4fjDt9F
49sfY7dFvGIogEHzo/JrRJEgdfLPdIeGR+2lEPXz8D+zpIOWKV+Zl5ciTiir1hqUfTRwftBSh6/f
hWNMrkCyF5OnfyrzM4vk4m6Dls1QZxVVUbYgVbrFEfILECIGH2A5JIUebCrjbhYCgWm53n3CK2Po
3Svz0/OJ7UKcRI/9vj7jkvmQI6AUUDbIfvzkpblHIILtd4QqJ3rOFbmmtAGl/kCxTYhcf8Y5QrWM
FxJOAfT17wdeb5EXJ6mF/PKgsbQbikSVtXGLiKCGw7ft98/h9msJdfD5P5anlT6mEw0RP3sFs8lP
DhO0fOo0IXJ6bOAZb8e1FEgSDgMpW2CPW69d32xOdY5LSBC0NEMgynY+8W2dwiUbpgxD+TH98jtN
nZkfwwe+Yoe+rfYr4NQca+QlurK9q9jaINdC1s9MgvWfU1az66zu/LgKZoo6552UtmV8/3rhXapD
dpEB9RcG6qde+7Iwj1DE5dEnrd1a76ac8pYLvfsJ6biW5hkubePSY/gkd4d1sXAgJ2+kfi6XKL3n
Djqp9vi5y4vIrWA7ynk+7URPIXAELUMB9ZL/AFkbV9fHjoPqDjxYCQLCnEZxeOoZfF4cdq3R9aQi
7ko6vpM7qnusH++E9Q9cqBSxTKt3yXYPcasyplD13YKsdfNZA154RsdxATiuu1ELDugpHCFmLnkr
HW9kVNGYdvuSa/dRZBkmWjgvUh9vQbI61Atbvn1dmCiOfLLq27FKaMSyEiRJCe1FmVzwIAe/VE3O
c9sfVlk0AEwz1aoRhv3jETj31ovHppsCPeUihbLt2uwyb7l8jPn3di5Y1ed0VOIH2RqRW1bNdqRW
37y2Nr2lnIujMnuPf+PKiPaL/GThqc0Fd7gyiYFVLtkiA7paRwofO2VS6pjIDQv2M7q6hpmtqTPC
2mKZPrRVD+IadJgj/AHC6B9HfxQNRAR1WxAOngJ4qCgIbPokOTHVbG/AuQu7x3w1RX7+YrgFV13n
gfvIHP09Wz3eJsXLDjOFKgiGQK7xtz5UAOusjTK2Fw8+6Ax3aWB8huiqcFc+kVfwan+uTroay22K
eEeOBchIsZA+OQcFq4wS9FjeLpttQAKf6OhZN/9roOeryLaLFU5o2KnfHBWjJd2CmTgWnFyzBzo3
y/qrmPE6qxhiN/VX3hXUvEsXqy2ldDXWxAWbhycnaSZ/NJOUTqJahkgyqI0RpmBa1nLw4KAiANYL
xdT3qlAHh8ruZgXRvte6xCmkTwVh2AcipKdHbs5D4ta5RYWFt2PxPSBrFaS76GP7sUW5x/cXn46D
SA3PoXnKdF9rkRdBGzaB0SLKuYAlEGSJ/q2ERz9HvKTHThzEuVjab8t+PvN4yDDXRf2YZafdZURP
SwJzhyy5QK1eUlYb5zhTStoNhlrX4z7PYvpZTcfK9SIsSqFVG2D8UYM9JZoNYi6B14SCr5rpWRnG
iWrTKbKFwbvrGJLlOrCnPPYEiL2nGtwY+U6CB4v8e2OOqREgShGgkF6oBR/4A5ozuNlWQ6ugFydq
P/EUqB3jBwOn/5V8N9nLnQHkeBZmyvwOlFkCDgoPp0OtuqxXjwBEAV/VDdAi8XJEmPhrn4r5CdTl
3EPrm7dz6Vv3/+wT8gUFpBcrZChV2WWlkElimVs6IA73oWK9IYV7bdRT7dc1v19TcIzuAgz2gWYp
EuI2k+OCxPkvwYH8j8TWa98En6T/NupPTI3Evrj9KGlvha2EEZlHOPGp/Q1hk5STHlrBvFANChxM
KJhnHlrmtG3kLZEn3PZ9W7aXThdx52yPttgIaiaEsm8M0Ac1oUrxLkeQuZTk6vsKr3lPPRIJwAAs
6gJYqUBa/e2IrK3cHa0HGzK6vUnsQKtQId15i+APQ9elLU7dpHwP9EcFwGlfwR/1fUDvn+xUUCiM
lJ+bhdSEGa9O7shVGAcuoxy9XKK3dZwkBA3alqmGBV5he2W+GolEE+Nw9bSrsOkYlpIvOaDad9wC
C71IEYgOmcIqWsl1WTc1BAHPFbZ0sfUcEkn5wyRMaiVfzdGkxT8IPpkzF+J/PAnBdWMxZbvFcEkj
MOC1NtJwUjcjdDT1G7+T4T/27ZJ1gp09fVgjwHIA/oqJ2SiSvXFjLyATJllizhUwGtGTyS+wsjeI
9n2JBmOQ4wGXn5wg4Kb9jSw2XvEjeNpUvmG8WY46sfTxvL82Zpljr3x75OOf0ElEio3JPyoaifHx
Tf6SqCOgOz8BEY0YrT57yfVLLynudLv102rsfai7XT2vC3IW/DyDaFTKl/grPhYB4WvHnCHYa/8w
kQ/SOVc7CsGlwi24jTS1+IUX8qD5laXKm7P16iXHYk1YFNLcZF1VMjihvbUzB42pFOpkEabzt85k
WNxk5ZOKiwpun/61VZx7JqZ0BrBdAybrxHNsjhJ689aApjm3bx2/ad+jnKojrJx4rzDFylI61w8Z
KyKvUHXRWqDekPNE59iT6wevaGvGpQT3BAiUoRXkKp5MgRkJfJOhbiO9AD/vR2ZqS/OH2YCDsXUT
pZ4aBle5cRKtDb0GJSHgCYCFwmS9bSkIPk7P4K1/hE8mZBiEPrDQwitwo78c9+vDm/b/Wld+dutN
4gR/xtVcs/PXUfcY4icNkdCm6Z3/CBXVheqdskk9TH2PXl0g/ERY1noMnTC0nEC8h7DmDHRjZIBd
TXZuqKLfk+OyltvBVHPfqkVSfUyDSN2OtLmN+4ukad/V5T7KmQDF6dQy5q3GquL58jxID7kfSYOg
7D1pIDo9Rjk/9GWuuzv3u3/rsHHsDG4hvLFgNzTnopTn6uZ7hsyHvh/u1Fbgk+2rAyRhwqD1c1HX
K1Smu/DQ4gOV6ho/LZ/dZ7kntBE2c5+SeOs/jqlBc3SJKh1mJYYcMERLWDg5LF8PbEy3+V8vXCg5
gTtqHvgJ4i+mfLJqLv8MndusvWqx6HdB2slfEbf4iqeulkn63O7TAXlT8qS3OyGhu45jBsqtBtiF
NdRP48HK3+muD6Yn6BU8di/hq/ACNtHFnu7iPcOhTG6nCjLRqRYv1H7bSlujV7MHaToyNuU7YKUH
hpgmGGKQG+ARBu0QHgX2qG2uTREe78vi8OCQDFJtG5N9NbGE2Q3KxmqDe36UoCxZ8t3MKrHpzhpS
7Wad5WM/K00LlKmzryk1Ie+gz9m+kmt6vBfH5pP/hsUe1Ot6+939pP68YJ710z6Efk7XC+2zYo2p
i8g85RFVtPg+9UMK3UR+1UI6aCiXz1RTwMTgVrdSWI3GCKPpr3LWrSPdjZ2yN7mmBwbNYQuoMJzO
y7CQS7DokpwloY68AjStVa6db8/YflBR4mBlqAmJ1Vtr9Q7SMqVOI6dM0/GA8dkS0VLFBoOQsuYi
U6MK7LnUlA3mvUI5IqIpWKSDxhS5e5XsXbAMobcdBaUpMdm5GJnWEZOitBc5WTLkEk29HmjtCaLs
xn3g9nsk/JmSRCkoPN3YkvhpwQU+WBwF1E7xOrGpqSEKsWEgqU3Ep7XLAvwccEM1P501sjYsynWV
hH425Z11tzfuR3wB/7qhkzEjIkD6iyNbs7cxTo2P5lCwN13Op42/Xs5f8z015O+8FhENTEoeVYng
p0acl8n8ZU1GzSC+BBvz30ogivuAgL9VMYk94jzoj15LtFW4MrfqoBAykFjoKBFaCDxRAgX2ep+a
rg9RbFLPN4qn1EMLj5iKkf2kt8kzpdVoeu9UW99UjfvXLqFZk/HROxY4ussldNIJP9ymBLybfde3
ZP1nhT4u/alSYN5DALeFzNf7PPRwN4gPrkmGvg08WO0JsJrpyTu4SwMVTdSAoisl8VXCh83+36bp
joH1B9cIRe6uUUI3VbbhgdJyccmzEi5LaxOBJ/34cN2vIg0OoUWarGvnm8UHIRwbdVAhe/z0105p
vXpr/XBdJtrxzhhfYrOc0qXngdlHKFkXzU7ZLdG3tiFAhVY8FPHALr+PB8Z5ChWPJV4o/2jhGdt9
QbxICNPiH5Irlxlb5yl3FXLsMm6CIwxtzYRUEf4WP7hM9lyaAO1QzpznVYgxHYA2gDYnJNomUTXk
c6qjb0yd55IR3AIYj0Nek5rLHP6RWm2Ssq3738rvvfqzsC2vVfaDrKh27TrBfA+aAXxnl8cIOQKF
c1EpgZY87QRD/uSr8mV/43w4A6YW0EzZPM5PoGwjOPd4dK/ttPWhB/jQ7CswcNW6D9aUW6iSUlVe
PSe595T+NT1tHSF8Ac77iLRKJhryuV64EgHvegZ1lVXFzcCKnfsJaIvehPhqWLaIwQTrTbvr8uLs
/HSSnARfz2J+E26DvLYfMAnTX9RqWQhURfVFXEZZE9fAgO6Xi98De7qytfIF9UmezYdSS4ot7c71
MmCBIH6bEbzyyqx1stNTLS6M03L0Momnc/iXvEiMYIyOJUaM6mpbaSy1V5YT3yMmUPI+naaHWjNJ
ufMQzbG4pBTNXyBnt36EOzcqx+Nc2N849zWA6J3D/dq8BJ670MQz2HozId7YRBUhChrqrulPtfnm
omq/i+lQMOmxMm+D5VFBkzjNT1IWgO5KqNxvtEg80kurXvkIIV1eyQSFEy88VpayqnUDhzhOUoz2
JdjgUT+TtB1fHiTNuq6M3XnhAbA4Y2R/JM1YE3rg1qzR/7BW6ZliRV9lIdqTforWgZQ4VR5IAC2P
j1B9bw446o5lo7wZLiw1kUJnnHXsl1+YW+6X+rYqcdaBkUnO1IBqELHynbXIDRazUNDWM0bfIkFm
ZEv8HE9C2qRmqbDdePl6F895m3kqWxbrN3xRcog0X1WCaec7pscg2m/rH8uMVSFSmLgja9fB1axm
IncaiWLP9yB7MyUqkCFpwktfi/3Rmg+oyERWgp7/tsqMXaDHtZv3Kb3bmjRd1ftqOy3x78GNDmtC
LW+Zs0XKAdWgc7xhM1uu/llYcVwskxlhMUrmbBYJn1WrQ1tay0/Rm/rKsk4evU40RrmlHcEPJiAZ
2gmDXUYdtCM9RQUUeci9+PaCSj5vyno+XNAcD0YtxYkgPX22Ttcewqf+2vMBjrmtJli7VOxqTFRO
5OOgOGhmOX7uukVWpANi+l7ZltQs7PIyuLGsCneTw0phsgKjNNYnh8iuy3jsjwX9JEfmCPfnJQOW
nevZfGIrFVKW+h7227kZKgf+2bOc2oCPJ/Kcv1LdQnrkK5vQqLIV2Hj4U9gfPkdrb66YmzdiA5FJ
miWTvH9nGGlfMcmlp+h2L4Uoe2VJaBE+YAe4RE9D5ELjb4jCWwYQoj054QBAVb9jGsqiBVyUcLyQ
VnQePcUw5fXrvZt0Ck7TpN5tpwf0oCRTKV1Oog3mGMtQObLSQCD18dJyS8F3PxzKuCFdaE+yOrYo
JJnGlxIY1tmiBg3VIkGsTWvWOYXm9pE7bPwhVtZDtHNKBBtxIxN1oWwQMKxXIipf90dREzvo5dGJ
4bf4aOgtdE5jyUbfJnz8jYIo8lY2wivH3KWJDnC+av2Dhzuy+JN3NS3f4hgVRTfw6p1GBz9gR8yk
xH/viafdA3Z9N39hfGdfCA4cpKbp2VcDctslsGQ5kRsJwqaGH1KcQuF2kuoYw8BwSpPUhdynxgY0
LEbbR/+LgU7Yghk+6tiJ5GRaQAbQA9F53X9/MBEig2ITQngxgtzFhKixfEJKSQTAvW2uPurYbxql
XBr4EwUgqF2Y60k7BntgclE0+KT9ZsD/jNUtcc1SFt9jWXMPhuYMJM9AZcNepx8yu9F3ZuMolXdO
1l2D6sFFQdAW2NQKDq+l8JjSUNSq4hqvaI29IVzfxgNsnnFk2x2qP2ZqezlhB3XVauSUV4MEn85W
w7LchVttwX4mIyGMxhrKvmemlyfPPKNYQ+ShWfD0LG6EzcmWUAynSqElWjyVovXlLfI2gaQeN8r8
iE1LVw5NNtiAAWTW957rsv7vCuNCwCVmjH015E/oOUyVSJHMiaWhbD+MhMf+DAwe6sBO0a+5snm8
P5rANk1Zl58MOr2fkHoTsy1gt+dLdGGgEX4zKAMemffTObaFdzlq2patY6a7LAPoIjb5Ugg36UY8
PChD6VnNj0NBeAjbDr6Q9wDNYEXYpvhkmiYrtcg7DK+SqYoUzZbswIxacqkzhr+GnLD2JjDiemeJ
wvX94zBfgP3h20Y3HnUZ4KNRBssPiZ/vqvhlP4/vHBHng7lPnkZnNzx4OzeaeVKAhDgiLCEkLwdP
fxQdhzox+q6Ax2Feqj2Qw3PYVvKgE0HjV8KxuakN1fXVol+XHPP72Tp6uN0VgdJCvR6S4wi16vXV
h8ZwMU8S8BLUgJTqBU/L6Mo2VT1RD+qPigASWDBDmj0fr5WCt/eAgp3fyMnIahgZpe7q30e1B7mw
8K0LXJQTyOr6rciD+J5uk+4MTKI1gkJ5RGAQ30cypQGn3TZ66VB1PVbeNrveCa4VLh93xxVCc4Pn
y9qVzee1yoEZTp2pwRqPmpCtIJM71gz+fe5IRe1qJwYrYYcVz1HwFO/GnozH1hhtM2uB+DsLyFTm
CYnlQhg1NS13JCDzbQSKBpLk/7fa/dSifmb+pItxBBapDvyjndgor82PLsZcZfzWLwc+w/HJ1g5x
LLcrB+/xG8MvIlUV0eyzwCw8d7KN+K+CC0nDEj0yBRwcRaEdDnyXmIV8iHegg/9qnWIOc0bz50UR
fXVOvJ0esmY4FPeOLhy4WUy0PR5XHVM7u5FuPvNyabethu22C2rCvCalgmKlM8Dipm2/R2XjFnAb
IlaYCQzjt2L5FFkyYxb7u6VRmNhathf6H0/4P9rzoFCnr5Bc/qj3qxFrjnyva9z325iHnku2e3yl
MQAKXLzkZddBE1Aih3Blg/DIOMn/SyeAX2xR5n7f9zlpTbhFIoEv89NdXPOXHLnzIYLAGzn1GG7p
2R26HEg15Nz0WiZscSUPTRFZOBQq2hxj+qzugx7N6d/PWRynXSWP8Dv7AuwSrsuuFcP0UqxZY5B9
xVfvyyUSfn7fsVUIaX1ozp4Cs8fH00Bk6fdB2SuKspLmSteoG83auwgmhSmCqR3zz8egERuhB8SH
0eTgOxfCYglwdvJV7kseig6fYpH91xq90fiq6ILTf7faWm7DkGKjP/m2BPQmd1/Ilt4P/mx4mz7c
o6C/ao3TKRPQlI9K2gZrxZa4+MXXxc8I7X1Sj1AVXWu5IV3ooBfVW0bDcSHFBliN1dcbH4xDzWva
o+1XURYCp83lhDp3n5qicbA1Ck2aumi9gymxN1nEyQTTPtXg8b3LnVL+pFRjQsLl8LNpIdcYtL7X
yXjd+Tm4ggtJa+NrhBzYozumwHY6y+qkgJsTbfIkd77mI4g9mweZ0Q2WEtKkvHe3grFwAhvGImEi
X/FqXCYXNN70xjgW2omgKTm4doTVYs6GYteXpX9XhKYSpHMCkA/bcoAaQEEDzU11sX50fnfj+B1n
wd/xwjgDBbBDMxnC0bBSMsSzj0LKpMMZINQhOdCSjIXPxY6UU2a4gA0bhuvwwYJzxDlC898NYF03
aACbU+rDid+5RjtAuWO9wUdEjePBVUKyQ5QFbpYpFnUWMJtgb1hR77H1XhBj/W5UfLu5nL7t1nKc
jJDoY+i2QW7P6qowBsFgRVp14LeTxfQAJwP0N/+/lgjrlkPwxgxJvP9x1yN4EQ/Q82Av9GQmIqbt
Ab0/JTOHRkKo7+iFI+PVyj3B8mwpZSkPFiFnV3udzkE+goksmo0NlOrYTeqiNT9gr2/ziS+ls1qp
UTtU54+wMtnIhsS0QV9v757CZyPM6zFuy+H6b68i+oyJMeZptdc/hKL+2mZB+FF6t62eNKiMFJox
q9ayVSaJ+7IgeSYdNBF1p19nOiLmk6BqozALQzYPR9k1SAqrkV6z+7bV9RLQFpKrwnum2ZW/Q9U9
ir+ZcM0OU0qwmwoeziRsJi40UqJfMh+1tm+V2AVqqUibzRr+r5zcLwKn0F4Bon1o05+Dzpa1dFqj
4sdknc1xKO3Y9T30411RMHjpOl2jfcD1vJAB7+lS2eGi74NXneMHYQPQ0RHOn4Pl6YKRH/CyZrIR
LSR7Ii9CD20I2I41r0xUlUCIMqvdL3ojVLqcqjY5dFiewuybrut6xCvHXx9oqETOVyW+2aASWBtp
QZa2f4Y6xOXmvkgqM4R0ZMO9diPZyB3AVdF4MoaHvVtHtEBN3hPprVKNvc2bKE+GfB91oM1OSDmQ
dTFFIkRJTRXc/5Znyck9CyD+kl4ywZbDKHaiA9jGkNoZuI+pRRVQX6ohDxlgF9C17qXPjqcN7Tt3
iEundIWnilnahpmJFxF0o5CwTMweGxhwfuKodelvtbpA/CNAbL4gA4h67hBOLc1i0ajAUP+UBPxc
BF4NL6clByf4kUTohjlJgGt8GdDVWK+YDW6XLxWix6NYqygXNVZvc1xRVroVOYmHjdMKdh1freZV
9RcDmMwCQFiVsYmOkxSYqA0SWEC2TaPXPUIO+y7gFCvqcZKOn5abVF1JetemUJbK6Cs6SWMhKe+H
5B3oUY6rSGKdga+DSxgGXRX/jHSOIRi5edlaGAq6wKyKmzwdRfzADh+ErZmCjXteFQFuo3QmAqM+
BjRHQ75Fr23VkP3KeSagH66AVvvS1Y3oZYx23BlJpHN/IGVdeIS74f2/JNt8RaV3SqqbvBC73Vti
0U1RMF67UcWnH7OuxxV/DQJ3YYj1R+VlVzhnAzKJJRCpSPlq4Hd/iLwicSd0nd7SLy/46PccgyeH
3ZiXNMQLmGh1MzuIFJuQfDIr8bN2ykXdCq3mc/tzAVk/YITY7pBSlpcTTlxRpl6AOKG7ZR0ABdOk
crwOAZM0tZ6vB+y2fb52pGyc872kGQqYlhfB7EDlB3x4qqZ4NSnZhhfsCYhN77ZizrdyppV9Ps6T
8hV4DTALz3ALay/0PXKxPsj61GuPZ8kul5JlL+1dnutZr3Y9mSfa8VUcWH85uiqVFMHKtXVslidq
RHrN0UMNNurHODpeIrs5+oAxc7JkSyUxexpDfc3e8UJr1bfLsrMDDB8VvFqaHHhrAdlG/oGRNOkj
diO7pzb2mFiHN+rpxa/tuMqEJ+t8ofQlrqnvDQrqL8w9mn6SyVd5wQzHlH48zVwHSstd03hVPvRr
BsPkdq/y0AOgZV0TO19RIU5mWJkD4csN0Rsc2LJ+bgXOKn76gdh/xSmdF/J7d32uYa2bMNoCvt75
x8YZhCSKH4Ckedqxr/HEekkYv7mhM/xnTUxPDvDdLi3UuwixZBKy0/LKuMIa57jDy9fFi4FwiuYt
llAWiOupSAdbqJHhl53/jMMgbkqw+nUNPfEbMAm3xLHk6vEWiw2WBLhvpevurM6zmgGvDXbkZdZp
TD/WdXGv0fVr4t2oFXiciwZjDlfHA6ITIFKVOswswr81FVaiJiZJb7oYQi6Ez40AQ2HiZJAbJ7v9
akd2k8Jod9IyHzyVG1tFVcC3io6n4w0Kv5fXe7QBQsDdk+mxY18ydGtxgXgS3qC4Qb3ZQtAhn61i
UCnbR+ancFAtIPQI8MrDfNl9mgQavFVaz9FZeBDVCY5Vp/h3Ip4Rl1E9/1JMeIkdILL6R10V0wJq
Su898NFk9ZRAPe3VFKMSe445SKrH3DCPGXnmX0DGKmku652s21xgX0Hrs6LJLYg8IM8GpwLk04s1
CuBue5tiA0YIu+qcFDdcKKv+QlnU1B50cn2IvihTJiGw0/tFnjFcSZ4HVXqRz9Umjt3QI0zhrcF7
0yW3kkXcnY+1m2RYPfDZdrbyHSCHzmWH0fUBR/xntccQmyH057Ru78z5tWL6+mEMH4837r7aFSgV
JkJlUW/Lu4v2c6B++YYYzEoMuNCWpYa0bv9joEqOYwUs4mL0MgyuQUJSXQtvv7cn1u373R4vN/ey
XdJCUsvA4yBSOHtYeAzpdSm8naDhnGTp6tbbIMJNtacia57IXQ3AKEwQGXPaPU8QR141V99JnU8n
0UoRpZmPxqmOEXX7uWtmeCxZ+gXerBe0DwwVYcCTbFMLnV295YsiDgf80Xk8aSvHgF5YQekCY0Dv
T0t/IpIZOP3CMUc7X/23zWzpTOyt7Tg+ixsEe1CwVWLg12eDx7OD+tQhH4/nCBqulvHERWSlG8WZ
0BaA0upofjaDhiRtAJKHVdJJaP/sKReyJ54TA8jqcrviU1wD9drAWzfr8ghbN7Tpykm1AOc+OKDw
YaTOG8uc/1R0AgHrXw0s91o8t7cjXynOgnvMZZJiBDpnglsUxv9KczuwQpAZitYedWoA8IRmYKDj
wY0SrsNhLzFcqvlHd2qzvaGH9jZLyg2StbWu3RybkTXN5YDUAYxzx5AppWozkbHYjpnNM4VNcs6+
oaMpfn0JJZuGolzX17zEWB7II9YwF38cv22Ud+lKF3eS3NWzznwbAkecGFQ8dUDiOoQcQUo8Hou7
iSnsZgLEbXuhykJbRHU8QRn4bHG352mnEvgvf9lS6hgBGIsAx2iTf/6jU3icDG/7yPvc3GhNvBp7
92oPC4q9Fb8V2lX1Nwm3k3AcO4HvjOEWh1fNeWGr63aCW8ZhlpbUugYs6DsvRtdl/bbYRZVRq3Wy
plaLAl2V9riFqLvhhKw8KMwptmZvLTeTHN18zJrzPX8m5KQldluC1H0BOXaGRqxqt5mqE/cAUZyr
OVFtHVYhZKJ2Y7Qmk/hLqQSaO0VQ697ynt8MKxXsOjh4P2j1AK0dscc7wHwVUrAZOXXQvN3naaDw
ie85p+RW7Jqdo5pMXzFdM6/EUTj39kOUZs5NqlUnKn+H+gzmyBQ5gHtDBuJIuoGX1YHeHUgG6FYK
cxvSXKHJOIomA7fn66wS++K0So/c8ClRLAeJjs5fJ1wEQ7ixHR4moElaooiE2H135CCdoTo6GlYn
rQyHCTHP0p0lJL07PLJWTPz7L7YSv3wWkuTNggjGDkIlhrCZXYCcLzufO7cfPZQThJzXyivQ1PzL
6ocy0VzmYEaB2fRphMhQXd+66mKETX+MX2KPGm1IbRXNDVW95iRkuS0ykQ+tFel6uCFXsnlqzoEZ
9KQab8UIeBGrOat2KvHCsWG8224du/CN/a/iQ8Ug9kWjOyMpc9MINr9MJ9zCrU4wnfKqhI05hUir
bLEiQkhcf+cxPQXnyj+ZK0hV2EdaTiY39j237DbXbNpVsU218g20HPYm4YKkgz9C7vFT3DQ6918/
4qMwWWlhtV+3Xxf8mnHo+tNnouv6q5Vy4hDdQmwF38ZIQ5yedOUpTUMbHZuWHzOhjuq1WkDlmODv
tggJ+bZF4haFy1bAMx2n/qCFf+PDCC00nw8Y4fR3J9KGo5yr3YQsm2wJB57hvWDpO2NvNQC4ZY5p
wZzJ9E64jg875kzJbSRyS83goKQT/b7IqDwmZ1GGA/80fdpPYEMlLC7k+EYQgSskto9U3aCYDHae
ioavo5ZUf67wM9fjjAPrNN1q5WboBu4IRFtngfQV0306xYxRYgqsOKqumGzUQ11A7zwmDORWflWG
E51cFwtB/1z9GUOdOzgBO6uFy5MEpKmzNvfFp2nBrDxrT7Jw4tPvaOpZZtW4wIbNXDRwn2WoxrHh
sTki2YiAEYELlenKNL68RV2WrXJvf0njlca3CidwSTc6HOCVNdisKfm6HRP8dCc01/vI6YrrOl/q
v2kz+cbfEsYiMv8Niva0VbDhu5EkBd5xlr9NFdFtX/GdvPrIGOJl9065fQvf/vBuTGMphxaA6nd5
N9gliWDDO83wvLQ99NfVfqf0bH8Lfc+MxspgZoDrHovDyvJs7ysOkYxbt4Nt8FsFZ6fQ/DEh80ys
KeCQ6nViw+wJiV77fh2t1hRwCnlEw9zEAEM2upagJJQPyMBMQHivJBLnzxM7U0Y7EuPXNJFOG6pV
wrZvV6vxqMYC6qU73+73fBIZIGEVrwEL95NN+puaz1yRhQdiHpse06bNRf0YiBI7z7jiGJkY18pq
7eolp/2acs7k2YLMfHgFOZLTYNbz8BCFbKaD3p109+DTgdS8H68YTTYoQa+4uSsVGI94+2g2BTLO
vyFxlTN+vzcTZaS+/c3GzsjY/SA62GwaeiRYLLcfkzKqF/W9IFEHZ71JXy7VQ//1oev9S/VQOJL/
BZ1xF7bPNwfE28OkUPOXRdE1z9AWe0xf5rXXA28R4GMWJCkuMsl5OUDm1N5qF4I9cPoIu7e/7Dnv
Sv82Fv3xdd3Q4n/RKVNZAAjjaDjRt67HAiaTvPYz/cZfg2JI+5opZC8uSLAKJ4wSZTCblR5JJt8X
YcjbAu2IvfVb2CSw9lA5+nHfhvh1b2mUWW9KXTp04q0DYhdumi3k+2BS/uwy/el5jFzZbA0vyEah
WFkIbBp+afOBq6uIiwd53I5KXctOFnTbGmIPKiux83TM2CYirjzLCbG7o7YoisXd1uAvC55kGokp
uK4fBhhs4bJqAqDufdRswL9ej5kUUZgfJ6i3GagRADhXzCeDpKgw/6n7AQpRUDBcpRgvyhIyJQtp
CoECmAAyCvp31VRxNl8o39DUPkSE9gBIADBEDmEb0tRgs1hbazDZD0LCagZpvgWo2nU6vNW9EbC8
RZc64XUcfEUQQaMH5MRDONH87vxtAO1YkmvFH3az0IEpaBeJ8RU7i0BRfsyM7JCO2tSPVUUJYmA+
LjOW0ltPJiXBcwJQFeB1xumu9Ab9r2YnW1sn2S/sN7ojsFJTM84rcL4bD8g1AJMKKR5gsg7aW/mP
JTQyGzpENIxvlsGwIydGujl8KUuwSMoK2AkTEqb6g9dBCrWBo9ryA3JU8VpZf5wYxEocb7WoVNdD
bqC7/BqLXLZiSz6Yhqkjcg2vbJA4q4BYmF1IMQxIUYpMKHB8blH/iqLL8PUU0z2KhaZ97/UE01H5
oSHhxZ8k94f4W/5wTonNhzb9QkLu66ScGrdVu6yMW4r+k4127hcJDWa1uPMm9Dmej7DgVHG5DdTw
2hMfbzRR4fysZ9P+faTd12nPcjTelv5mmQSw2SyzUZAAFbzo+PHtZuvC6MfX5f7v4PQA7lwCUb/C
7r6hWN/zJpqXDW8oairOvMHKqro2ZfS1dHCog2JcQFKYyrBsiExWO2tWxQ4eqv0cverklSp4DvXl
Gp/mAFpjgzNRomJ4q5wqzEWMywtrc3Mq+Qcbrmzn768dEvqSMwp0Edz0HfYdXNjYZdcvlOnNBu+B
zQpcdJ6NrBT6cpkuSx6t1Uk8MbN+A2DRWxnVSTt8YUMdE0rR0Hl4X6p6534rgPbqpKA2sYKktWeT
4pU/HKkJC6gjArGO90tLZKG1FYpqUXq7gkp+FevsBjeTHPgYqHjHruKQl9PaYNgEQk1E1E6e84+K
iJ7eAlV52mMYMJC6lJ6d2qQmbAE7Err6e6lkUFgrHxkJ6Iu02y3laHQ8y1kQM/i7gZcBt5VFmI1N
9hpVnCODnlZDuqjuf7lyXeYN0QlSjdTS/S++Hmn/9IzrgjwhfXHLCfUutO/4Uqt0m+KeZtyHDiU+
NHqJxZ5i4yQs3KMjj4cGgVFoDpyzAXrNtxYMO9S09/Y24m0nmcEBkDmfnQgPDG7RGLN6uAY4WqGC
g/9l2W1ckgOQRwRCsnh5+4IiBZvr222njxkUPyKNsjUkOM+INsTb4cz0VDSzfdxGRoSZwYijOU2P
fagT7tFFd5uULuocx/DdHkykqZUzh25A6ksAHn/BLfBpudFgpbwm8I6qeQy4rncWgwQlrNV1L9wc
7i2/5inSCwYA6dRXBvb+EiazlJoh1djaml/dZItrGyguiS0Ak7/DVx+4LaJNe/ZXriw7PHXs6Jh4
m5sRdVW5G/jPi1SONzijc6q85dzKMKxCsRZw64nb2cGFy4tGfaZEq2aTgBHlw2broJprqgkNKjyS
b5ziAZK2hqauE2stm/LZiAKrfS6FLb/oNdR/I8JT8G8XV1DKgIvVaIAicEm4EUX0OieEUin8WcZs
c55v1857HCuRuSY4kL5p7FkYBrbZnIqfhvHd8nhfvYKbV8hAaZZQ7uwkMMSfhTfQS2rcy608OrNj
srPWiUtC9OoMGAfsIhks5MAhDp3toU1E+BAQtAgidYu18jA5NYHQ2GvVKhqT5iZKjZBEDWBd+4LT
TMiKsH8xsJAPR75yLdmJR39to4gVTn0Rp7htuVMFyBjWuLTK5Y/OE5s75x2m6Chbwk5mSPzVf4K9
vy6NNtKECnwrZEotE6CZ+hTn/XEVWa2T9p9OQ36GK5krcuHNmzKIbDs1UVgp/PVVzUpALbGdHnAr
mlWuWkLGBmWJs8knS7WDJQ3eLSNEOxFlCmnhV1vSRAtBGVQ9X42pjrWSE7vHtni0i6NNtHcoYyKS
JX5I3az8kEgstk/M9OWQrSRyaO53j8LBYRYu8xBrCXTxJKCwSAyKwgAHvdqCBn6FLVx+KX4pg2bL
58K93P90cZ5NQUKCW17SAVfqvvgpnb93vpL3WYVWj+5hzedQRN3+xztrmhWZVXNhh9Tx8h7zHnzZ
5qbMK5qoQ6WXcgdT4JelQ7aKJsDuT2VgRR0cRGF2tAjAAW3bo4dkMgAWQO+qRTn0C1fYz3IpYYLw
SWnfp2NxUJyx0gBm3eXl2wLkg7tO0aJD6FowtF3GnbGOpyHhQeZ1fqmPC0sV/W87VYKZ7VjVuT9P
XN9RDtWqLSb7T6bEXjKEctsvldhmKV6oNIKbvNxScDW2vhzesvzULYAJgE3/ieGZNyzIHRI144J1
O+j+7wHlhxWVP4i87C4qR0kr/mOFXfqR+783lZ9N//VN+JX+AF9axepHytHBINbdVsOYD2vCWcsA
TREIFA2PqtwtFrScCFESOZqAHK2TlA6Opo0Nu1tQMRyhEwO2duo6ppCaglpvwOY20v4GXA05XESt
or/rfkJRs0maGowHGORxNxp75nG3+vyKhnrDnKeBVryRknHYmMauSw5psMWfKIh/QalaPE6dfSDH
E8eiyVQoq0cg3W41rrdBLf9EFi+x2nVCvpCONPvRceBjei8NGCZ4gwt3yrRT1lrgJhLngCNQ9h3w
UMSTwS4+SCm2c3RA0AB3G1yKhW5E85orJOGWZjfnGrsWgCdRhg3yydRRPWBnbo0cjew5B3PMM9vW
duIpHSzpqXBMi5MZq1N0UBz7/+rMEtuvg+EGW4wRrB3jjMfr2n7bADqRfgkSikCzewgpfUSXFRco
V6fACNB2BG8EQC0YbIwtyIyyK2JGN/BbJjnqTasXlwNq1NPYFKQvOtQWTiYcoItngINYYLmTWIzT
Ifmi14amigQk0x5d8iyN9VirBglHWn0SiL52eRnz+3694PU9f42Z3VR3omljxI/2CJ5XEOztbW4h
t1EDHH00o23VBWnrjPUHcB4K4bxk3n8kbPjLXoHuhGsmHGQ73wyrvb136xec0pFSROM3mnbCr54O
zdc5KnfBxqKXPrBh/xU+1FDb7oHdvTUvCWfIak47FkbmuSghgOLhdIOK3eY9ofli/4/UcK0gigvX
3V4uoBzNGZUcfGqe2q171rUJ0G6kDuZens0iAg7IKUwkhIfx7gG4VhDOi9wcvrwL3p99mTbc3DNH
DayuliMsNM/1nCJQPN6UnDIwluCtkYKQQ6IoGZN7REU04Hcocb6YTtBx45HBIKVk0suozNMLe4wj
2IoHkKMvbHxrO+I8BNrsZKt+P8Q4sYhFXZ1TcuxrnsW3eqT08x0NTLti5UE1JEGjVJml3s1b94R4
DeGFG0cT2Xq3Nx8hIJNk+3fVDCU6QDVcykXKDUfn5/GH8RX3Z87rxOLA3NUiRS5AJXHTdT6sM/35
G9seyrEPVKnJKURukiUUaNVu73IViyFrBa2TpETmlySSI8VNBjcJQ8k8jourtVaBsrnU/Dr9aQ/f
jr24Sl8eQ3P3tubY+CSzMCh+5OK9aHxGpq+jAJCiDa72Djk/Euy95DFi5Me8aP2rMIYMXctYfI8F
Hn+PgzP8UwzLpynbAta+5YnmC39W214n1z36Uof/05c0Kk4x5u3oVc9+7VIF9PBV4bNbDrAC+tNo
Z6nQkXG2m1iZDb3Gw3mmmoD9tlZyhGlLmxAhZKO3thKqOCwruUDyvcXcB+XYuSBQOf1oaBbphgq2
krVA5W1kwkkFKVHJnvoPZD0X+ZiMMoAAquK4m7nNyDpRu0j8OkYWOPN8LRosVhm9Vip4gKTw0HBr
s272WCKjcZMHvlNYZZdMfm6YoIG3FUqx61I5/ZjEkYXBgU+yzYGNRixuRj1cg7KXiuEU8k7kPMdP
X8TTB3PW5AgNTAGFfpDx3t6SjfzElTrqVAs13x0ARkVtcM1Wwt1vxHyZQybqiWlPReTvHEwIoNyN
JsybBaHD0QxHoWRHPaqGXVC+orh63I8SqZXUQxeSG/fjj01xZSNBVOLZaTX9wXZ3M9nmb3B8JEqO
cca9/JEPF33nk7i0/SLQ4sNL9rvFIj63MGHrgBZtEcg7vRrRpUWSy7s7rqBPKLVlVvpGHeQALdw6
wCDOOd02pHEGpN/NTnzSsdiJCj4edjmEk6T/hOi8TGDop3iXhhIlOJ3wzBVzQ/rR2jBBTCGAaKBe
jhc5WO6t44xWL97oU3CGpC9vdE0NY5ZVMJavDN9VRYVNE5MnB/arrrDvCfOl09BcQDFV0TdH7XyP
+DzpBy/7ExrwsVkr9agl/isi9HsGIwOKgO+T712HCIlUOsHv72exEw19J4eJu1POR33H8FHu9BWn
DbY8TX/3mVk2KCQ/HeeqPmgkDnjNZTKl1in/ZhVyZFBvifztEOJdaA+HwlnzJgaGV832GgZRCkLg
Qs88dN9Tkca9CtS7ywUY5EFIeemNMewAd/14qBgzPIcGn+GjmYyl+oWs35gWNkuYLvtKJ2zmvKs1
uqF/fayThUsSvoGfsUgzpR/5BT+PCRc2Zjj8C4EEQhOM/w/dTAXr9AHMnfb+Eg5ZYmIXqTbkuZKA
Go6Z6ttRTMf+uuKdBX5qIyIFuwhgrFvolCPZBtuXhaNqMHgDOdiCn4RWvAyn2V9Y6tG+RVypWYaw
x3CMKYaAqlU5zDd+EkX0C7xo/EPFE8p+kBnRCmdu3yX8i/ErofAo/ivLZfkIlIy5a5zoj5KfXeLa
7+thM+1Ff+hIZDHZmF9nJHufgdL7zrsLYf/wYumxJEmT3T1M0MlswBzIqtGv9ZV8IT4DYQMRGiXh
J6PXFavp4zIfDLLvsA4nhXDJce+wBq/fw6gPwiNvQNRVQy/dv1TsPdLTKoVQ/8MxGCA1t4aa4qM+
bKktSStav6JzLT2NLr4ZTV/F7Mit2+GRbc61tHBXCTE0LMg4w8nmzHIf7z1JQj/HoF89r4fFO8Af
hg4VhBkqJe/O+ikTIUn1MYD8dcdQEdXRcOTQOuBfZR/pl6d2zp3e5wFcAgd3pAZburqaEncYbm3N
6YelZqXz1o5WYdFM+AgmipoDzq/iKnoL9iIriJKSEiaJNIKAyaxw5vMCPMhEh/az+4xO/jRMv+vd
8Yhklpn29oyBeRwnrQ6C0YnFQtVs8GVQuQsPE0CHGc8JqhS9zKafOWAYheVOrJ3TRTdERIqChiO9
naj/Lq1BlKUPd8+QAxEg5pUsoe0TWhSpZJbhgNq0wVAKq2dCw4DbJ5MboBzwx1HYYHqiXjbSbCH1
DaF5PnMUCqA6NJDBN55yo0TmH99RCSyhUhVTG+2o5X+EFsKYN2OMYJLb/k6EUGMNtU3c8rNty0Zh
HHCM0LLJvY/LhkD0vcotkIyrOwtBCc3gd10+ZNoCG7AFa+PTuEERkwAEA3okj2RGY/CUN8myrpoB
BRALv84IDCWscTkq46/ditk48PHQrk3otXgZmG7+9EFYZJf97GEHYxMPWuzUSzVhK0RQQ/hcFJTK
Kp9NluL2d2qBeSyiJdzb8K3bQQ+wcFm+gKFsm8iepzKaUiPhZm1YZZLulTHgEHg06ElKiOuE4ULB
Je4toxcxgPutstqmpy6nr1M0JmJCXDq2XdFG0kiOaqkSRWnBNQJLgCbXsPLY2KOJstpi6uLpolDb
tKiYRC/tQfZBa7RvcMZ6pXNhdQbCvVBvzS430oS/ZEFdJazyrDnSJfn2WUvgfOcFv2T1AVGljkp2
nUGiOOSuEYG12HZQE75HZirpvULnFb23TIq07ey4I/MEFQ7qTH+Hc64xbNF5j7V6mwTkasBlcKSp
Jr24zS2R47Trn6nwY+L2IGRKIGJQwNQNe2O+O4p2FIjT6ZpioBg35nNm5YuW/1ODYWUNvk/AbXrP
b2/hv57Ti2/QIIDpCOjRN5cnBUL3MJJdwSHkUO+aiXuW69MSAEsCgWNVr7Btw52StZmX6P++JPKA
sWb16z2Gk+z4z+/zvUx6tOd7Knwo4VI+R30AKj8TPio5DpaVdvlerB7eDpLEBqJoVBsugVHIdOIx
Skhrizr34Pl6U/keXmKbnFYsA9uTUK2stSfkndAS73L1lV4nvprHehrPexrlGWnXpKjgxVZwEdI6
2105U+iYYhmXdxGOrUjEnR41twQWXwkDpWybhVNpcTuml8WD5T9VdF+OTK/kPn+DJUfrLOsg+MIf
pK6Z40iULykTGI50dQ9Tct4urfitt00DKR9wm5bkjj+Ax7i0R5UU2UgOh277xGQ9FdvcC3KRhAtU
TvTEz38O+dSoLGgndXmYNHAOdHWH7FX4/iLvHNwo1ZUt74UAAlv+wJkFyDveD17bbdwDygFeCajH
bVU6xsa1M30CY4sJoWAlJ6QZcTQOXHrUlk5NuHXWVDIMragWWCjqs/AgejlL0OMqPtb4gUzGuHd0
mHle6QQ3dD1NM82TO+9mq5eQH7Pfmo1rr3VBgb0/Ct8G6rGqlsSIxFv5mbNTT+ojGQznuG71ntk4
i2VJREnd1ZR4qgIBY7R4EIX5Az4ubs8x82ljpEltNzc1KDBK1K1vIhiWN20UmuXrxW0weAKub06z
lNc9NdU3TCAhJlMKukIj812YixIIeQu8u9AqgAJEcL16pZ0KWJ2PSE93Ljkej6GmoB9HyzS8a8Fj
SgsQinzkLn0WXeMf5LsU3TsXWyVR0gY90h1+AivqNvJiZDb1waTo0iiFGgwuc5T7OijML6Xm0p4/
xo50Acr0cJ4VTwG3PdkenTYKl//Z6h4rDLrnsQXkLoSVq5ku6NB1cOM5Ay8fDzp2NF3cDFlBUNLl
97mKtY+5FG6CnDQf7VxUabfS5b3faE98CMJjUH9CoY6o5QLLvAL89/dSdL4iLpK7ehcGdxfLIlSN
hXGdEIxaGkbHUsSEHNUu/OZHmObecNThX9o/4PQh+hftEaAq/g5wy2bhmr0oG2YHaK9SZrnCnF0c
HOGCVKAeZCxxmJRTHcc2DM9ZkMdYpg025PKsCKXZzdaGOaNzOdnYdipRME6buK3z9mX2ArBPJyPF
995/16OP4xmWzB8WFKqW7BNijfCvRQP+w4DubTx1pEm5Lp0s18iN72ImI3NwGIqWGcLTapNo383W
W36bxt7o+oKgAi4eYrgcv/0cyuuzk20/JE7RtZAG9b87e6tE2CNhHRBDS9n54/Sr40NKd80bP4Og
584HYVHyWh7jTSNaF2WJcpCALDLM2s8p6TdKqJTMfo49k1xOQnZRwzRsJoEJXdw31frHvEzqbHJl
gbEk6atTh5xPi8QKzaZqqSWxU0sBejw6EDHPJsGU818GBd238UFgk4coYn+0u2Sq/2Dj4aQHFrQK
tudMcoU/ldfGfG0Y2NSLYsvSlgSE4HWKmhACFvpCHMVmyx71+4+NXS2/96gnejIpMBFUowgp5yYq
hWmB1cDRR8RGShChqVOs6CkBKR2b12K9EjeFZ5EnpFQtlB8gvU+9cKMGET6LJxFdrJVZaY3Eex8K
qDCHhY46rBuu6n/Wcdhm4bpvDJCwLpnxRce/fwfqlLN8x6+okJd+KipthzEZo/3Xdf0SkWkhHepU
3GkT1wugvfavfrr1zigbJpvIlakak06Zwas3BeXL+WjLgbBKLsDFP8LyRxXQytRrsVted1Zjdwor
9yzsPQAaqEkict63ycAKetJqu2bjYoJVHCVBQKk+jKcSIZXFRGAx+c3pju5tfqYtjUb9kuqoR9Ke
G7TxL8Ciq3S5KRpEO3fypypRqij1di/TgmwWS0YTd4Ca/D6MMShovlAsV7125Dr6vUJAm80wRLnv
DpWF5eEcbr11sILPtUH6uHdAv6ITdci/4EDBy6q+9eR7ZSYcu50IWuLsFUZ/+jeFpQ+333QthWG/
G5JPjdBAhhexA/r97El6zy+unABApaZ3c0ICjXXxZx37JA+AYjjoeEddhuY+6oF6VGlANq1jT24+
UpMC0Fi/qV+TSpv8FlE2ip6IaP0n1ayC4DKvTOKRaCVeOP5z2pGZY5wLJu25qutDLA48dK9HTXv0
bE8ljawbjw1hUyoQ4CbbL5X+LYMEq5tLpcHwzdaIQ8EcMjYPkUZW/8fpLufZWazhaTYD6sKgTbwL
M1rx+e7wY1wv4IGaDAFNLkMDiyI57asoRi7W1xHqTbI3rpi16MOCAdoSe1p+e1DMcMiw63JSNnJu
AqcRnFpOvbfUgrAHn8vlprZ1m/DRCbcQZ4inOPAJjhuzu3jgyK2PL5nLddnCOaostJOWUmVG4ORI
USUA/QupkkGExQGietxuVaE6V8UjH2dQLf6r/+AXQOp0pZjFh5GDTvXemQmd7oRFxcRjhr9DwxcP
LJa+LWRa3hQhr5In9WOyZ55TRVR0PlTzuO8/AP0bWlxwsgGY+h04GOwVbT7LW1+foisGzrMUzlma
SMJq5urnl900m89NGoZnvVKABkeGG9gdwMiItWGDkDcAQFWtN9sFmf9gOYyRq+5xTlOi+K97VkEv
gtrNiMGs3l2M86Bi1nhn+nuQxNXwgug8uvb2G6yUY/ixUMAtEmwoMfxJsadmjQwnlkyJfj/YkaPa
mPZMCQSnNmrMtWKKam/FU+DxrTZKbJyiRxofaDIVid/+rq6riADltLLJmZo5pSoKA18SFDJL0PwT
tFAn5xxTU7bqEoughjXpTNASmp03No6Cwt/0TD/eRFuWRNbTVbJaZIOLePCHhBzgA1c4BhOXb3Pm
gz80c0D4fa1cnkBCJo7YjdI+6qa6IGYI8fcVHy21sLConVWk8oxeE6kSQPYGyrIjHhEoGgKxR8f3
efDAmwlzlSZot9x+E/740TOGWu5stIyLrGas/0HUR8VPe4317I3IciDgAMGaHYut5stFsVLsREDS
faS75EDk/oELFjStTrC3Z6nz6PdjVC5lv/Y0hOUjWzu17AHBDC9l+HeOoGQ6JdMONj1OOoDTmnQT
foDAWkL5muZO28w9tAc57K9thpKGZtOzMAwZ8F/Djh2QFupDR8OSY3OIj0VqrsWph9FhTK3Z23Sm
VBXpJ4MCSZL6oGwQAMm191cGj7xoLszl9k6nMDGXMEVrTX6HybU/odQAwMVRyRyUjW2LPeKZKAAa
fP1OHIVOnw4dN1kFiFj5nTPyQ8bCK/33kCuD/4I0ISYOckkH6W7o+QRwBVpVGtT2lbQKSaJ9gMaj
WNTKgpXZg1SJUFsTD138hgGJ58XDZ9R5Myfs4YLWcKiGVvZYU2A0MBZsfJ+CQbBnPHDsv6siB1Sv
Yu4LNaqomkks6sHXR2gaXVQKSN/DXAFMyU+7PKeIsGZT8WuwewYCQDapJzGjnjBl66Z0Nkt5Exlb
j3cixsyQkKHQmcgG4J0lQlMqSYYUtl6Q+Jk+6TKTlVw7i1v3EZGU2s8/cO3JO5oEATeCSLG6C2l3
6gRK9dARG+OycxfXTruoLGqM9c5NvjFgglFvBem1JesZy2x3Cixl3wdxQgFAlKjZZ1oZ7Ad+yFV8
rZ1QU6JcTqFrWt4yAE60j3HHBQf5uG4IYB3Wvj2/SK9GFFo8eoHGgEMCoVZGc64YC72r7cZBgNg9
C5y9V+cgo3L2ThtfMCxzLbg3PI2TVkoZWLQHR45TD/a9abRN44V5W3ly6hbrOkGYOenSNvVyOCht
9v/OkDS9jfdQ80SVWFbSmVOpx1ULPDFkhC7WGRzZ9/tmUjkKgX+TlihE19Z3ee7OlcuvhYbSMdu+
J36LctW0fSoqCrRXsGIYLiGPpxTtMwDiDuA3KdwEZxkFouzvDbiboCT0RxnPcSKwP8m+3iHgb2a4
j8Y+eE5vxVGahTAR49Yqwo+2MpfIHZaXsWmO+fAUN6Rv4iodqLKRQnLagt+eGnIPqT9B86eoEHfi
dQwL6IKaX2vHOgbRE0QuXJahtk1SyhADAteAjqcgMumhVg5phSomKUuHGfMZxP0MHr4KrJuTxOM9
Dgoxhl5fIHT6UcytGQLVUXxGIXwXXrZN61+Ml5GyeothFAelt+y3BaVcluxq6lPRsKqDpZ5LV2Ac
aFMGan8bJL8OZMEMfMVGC+hIa0RKrwiToCqBElgdepKYgNZWKdk/Z22H6Thnz16GlHqnwEdKEjZo
xQiUWwUoAtPbMp6C4ce7z2ChXPL35sEWmBZSF9NswwvCqysJc1kDa98VkvFM8Vuka2kws6YUKAxE
5irVgNBfsMM+OABnvPqA8t8waCal+zFFAEG1kSQmhJkF5HMHQcNZY3g4NhTkgqu/UKtdrcVEBKud
wiJUHofQaaooKngoTjm+pY6UHgl52Na3GESJkokhTMqZQ697ajaQdOgsBwmGAkHgMxK4JhDagfPz
S54ceKD02K50VFqF02wjjkQuUhzWWYYQhW0bBd7pPMai0/Q+7FCp5foA+WD62v2d85/PuYy5y5uS
L/Q2C/ySA+mTKX3SgDIbjzkNBuyW05x5mXMbtnpBCmqtn62RgopVgElB/vNMLbgbuEpC0HKA950T
z3yaVkLLeXuOGbS4MwxjM0pItyYkzDg0IGtJ4oD2wNhRDwvpttO7PeUNxaAO96Cnl3YCkFzBxK1Y
uB5RXIEEXLcAYDW2KNn+jRSHGqwPD+1mYXiz1dPxSE9pK+cKwvV+OD5sr/CjYK4B+a65jWmib2QY
Wbe6w754mXMujRAd6bUaqRQcGx5wRrmVxsSYZ2TPWg8S53RmvpN3KDQ8mMYM26OWVW/zNY6jGzYw
JQ215nxOTIKWhMsbv5diZCQc48T6N/6fnXTIo6A1T6iW3cxPZpt0nsiHek4F5MID2sC7pmrn4nnE
eT+lf71z6I/AsWR91+BHkoEuP7DPSXPExUPwS3SXrOmmiIbMAc7TVC/F3ATbmaQrcDNe/ciWKdVZ
KMvTIP3Pdzj+LXvkcUIPVp+KOCpVwpG/w8qxBs3eexYUrrXLX78Tc5DvrVOFkOVwKf/Ld7YLVnAX
U0yswaVTQU/ups0ZBPDK0cUheFGClMj2mDP7Bl3O9hFjXtpivqoZ8DYTAFUu7Lieyj7WctEUDvik
hy90d1UPIQfWGRBYlqT4Olc7xeOnAoMXk8xaWvq48DPbPIwniW1NiJjHvS6Y/IwNOPTFvMi0ktCZ
2CEbwfnqXtMHNp/v1q4r/K/AMStHHxfZ8drJ4FdwAYlDCqwZj0QssuH2blFpU2RJJLrBDyC1pzaJ
us3+ZImiheOtvc78oRWu3rSHb6m0CgUr2XjlmjYAB2IB3Jy6nmm2tcP9pU2oe8H5ZsJthXETkcdE
ujlxB9chD0VzZTgg3SIU/BCGri1UGDJwF5NxeVmOZUkowDLsJnBEd7wFQq05A5WfZMzmjkYew6/A
SQHUGLRTFiHpY6ZGmhqFSGRHwv/6oRcqISCAS7bncW5a2cC4RjqjcyNDW+Su1+o2dpbqrEnBh4NB
skc2xx62BAF2LJV3oBJ+lrP8mOvDE3p0VUN+pzPJaweyfUf5h7MGSm+PCJ4OsCvdwJlRGXcONZRR
CjZke0/asucwOmGiWsui1YA13ymxltCWvb7xWkMUELL0XzDcuWvPgepmHHcoRBynX+qudqHKn7+N
rTs9pcu1ouwqkeel8fspdIzL4I3SQjCjzZx/Xu54qJNlXOrX02rz5mhl+hTE5YXNkEH9XnYZvNXj
+yui+O+rdioehItpm4DkNrLzkQqC4+G3QV/J/QGlm7/1nyZq2mBQ/Uiu+Tk/yuUuhTaS75sHMF63
eOWPwVxvqrHE3JqWC49q6jKrt63OgUZbiYcrJ6NZ4g83X0NhtE7LEEj1GyPyCVkWnRHzGjxSm1Gs
iSY6SNLXWYS/3vMLGZmSCFOoIl7e4FV3DNqDk0V8tbiQxa95qflYtXaRx5Nt5lV5/QAXfh2dtMjX
Nta4ffMNeDc7tWBKCjtwNGYVigx/iPx69JZ4MJ+Le8dkPg05ra4FVoBbGtljMEFrhduQ3XXEddGR
8ToxYxw//c6C3WSvW1AWEZlocIoBNt1nblC8VQNvHW8Ynsf9xeWBiYFQ28bJmNoHm6s5fEPv43qp
xu42eJmFDGqe86o7UBLRfXWErYCVWp+7cG6G+agOmPUPpAUDVXjdPduiD/tOjIRCM8Y6aoZgOPa5
ohG+sSB/WA1CoQ1A66rFAJGRANYAIvb/Y4zrjl+LEE3V/bEYXXU3ffGwP8EkQge90SkxLJr7/B/x
O8Uhi/0RE3nrxQw5P6A1tASMXqbq0rZ4O3rcJzHcsMHy4kVqX+S3LLUkL7hVrgCxsCzu77jFqtom
TpPpLcWkjwEwodPy27qLNqNfTvjvRKEReFZm37K87SIw6CL027sKXrBTnx+bIwFUX69z86sWrskQ
LcQG3Wy3Ek0iJiWyyQ3lFSrIyecx8OSLQlM7GoxalVlvu+jd3DNqpZFBB3mL1g7lsRnCW+mKZePD
XzEvTh+JWMCQcr0ssKB0sGS5xy+SDPNbf1vbwiTAQzG8sAl2FlBUUhH4apM2eftJk9TfeMEDUKCi
I4tvWmUo9DcRaJOu+NSigINnhYSkQqX2GluzrzMf2lI3NBkjoTF3GzYqwhHcFgzRZox0gcii8LGT
eHKKPgv3NLkpPpnE+2XKwrOxXfTkT/Eu1BbHaljFZ9vhwH3U3E/wWubo53CsCSK0mQ3mr6pkRZBk
OeGZtj2oRq4Zhg6zOF337uRMigw6ORua+VewrZ/MG3dQHYOYQfQn672hnxlVSokWMZR+0r/qZEv9
32uk1xFzDp95tMJw75MOdHVKYuX3JOhJa7PeIM9VAWT3tWvBKOHvnTGEdMRefcWZO7WJypR3tlNO
Usy2wP0o+Jc4zFfdHIcPVSv544f4i9Lfvt8jfRSdY2MKKircsovOSWWb+OMyJBjNUWU5LOPxlDL2
EDX1VbLDhisLAg9tJoGFKlpW2CakqMA2iEv4soZJNsKb3MyqYcWGjBgJFc0aARjbf+1KU0+86L4F
8uI8TYFCqVZAi1NKsrqIYf5FCPwTuAlL4vySxTfNaDPFKhj4vVhx5QLYx743VIxcKabXQayB62LE
fy8F+MSUUPdQzA0kvEoD+x5yRrEViJdsl4WqGFb1OTtk4VJrYN/W0Sflbqd0kbR0hzLsS5eR6eod
oaM9h292oCgnzmLUfGNWuKTc/nyAr+FJI+AtpVtvKpXXUJReHEhOSpyxp2fQzniMLCztyHkPg5lV
smhGk8oMfYqC3OZTEnLpZ0uVkTEkWKmWTPp3M+5slsLxbE0J7YuMlUNzXCDHRh8OYy0wSxG5cZsz
X4914onUhOvmFUHjtrz0gxCIa+Fj72MqfZOzk57c16Xx2mQen+oyiE5xlcIALGFXs/pO41iLO8+C
RpwuKLRF4Yk1u1eE1BpipfbkadvHc60quXFww/Y60xfmhNQkrD2jhEw/46w+2JHsg/Eb8WGNYZUK
lA1Cdb74ahorP47GOHKz9Z1m7R1GzKXP4dZWl6BLhNKVez4Mw6twn41iseq5pCKD68XoLeleWRKo
mp671ds1GY2xEWjt30GCgpeiLAGRNDf/a4ajS+z0wCvSSLw0kWGUKbZq7mYbrl9tZ02X9M7u+7hQ
cf4I+668TwPeaxsCOi1irvConU6dSnNCgkQ8D15KyP0izPG9Sr/y6yYEAGkxm8661Qkn+c8fOu4h
IbE9YGceDGuti21tRxaM3WvRUGsW9anCIjlNo9kCpwOiBsH0UqKthXm5wKY1LlosHyWtl+2fDLtU
+kx9ZS7Fs8kpA5qT2UsxOZLB9dVGRoFOjrXqd8mMud2oWlZPI4iBmayoRS8nbvisU2ab1Xgpa+Dd
EBv8W9lxKO5q6pB5TN7hmwyWmNUmykr5vvBCGmlU3kif5zmZBot1i7wkePmH1EArwyY6ZFZ0tOY6
ISvfLnm6I+Cs6QvSv+6POPuXaoc4tjhwJGjbGwK5k/cpnulGcgiFjIXwBdhtWju7Xm+aGfNQclQf
t3k69M5Ru/nArEwBvBZaKYyLBv3yfyFqA04eqhrFapq2CrcpIBZpc8JcXjLnkgPnYDj/wPnxv6YW
iqNuPctsvJ+FTsk85ruTV6+ZgnORPwNy4kB5djtEBgWXD8tLsy9cN6WiEj9+EkxBWkx5aFWXnVLi
osw/xp+cuRZUT7AWuu5UTqc0wJrrQ/gmhiduL82/XgGZDKpCiN0h5URcVZSVoJT2lrK1pczHDkII
6w57nU148dwSDglF+10ImrNv1QiQ63ABgresf0IvGs0hocfnqlUUyyTvbzRKVnvhV06VIkub/+Aw
pHXWH4RPHhqCbzMLY2yGhJXiYjN5gcI/uN0UOS67WTjN5NFaPwzHLHOpWl1FN3SzPR/TuE6n9oZg
jMF3O3HTC/V9Zx4qTOoldW9pNbvnlH+iUtfhIZf9doZwTz5ikf/56FCUgcwOFWIblUgoDXjaRj5q
BuVZMwZxw77FYUi3PMM0yABIZdlY3YR96ORvxHb0SaW2HPZ8nfoBru/qOKgGLoxrh7MidovTXEDl
fI+Yh97YFyWdVtDOvnFx/dL/217Z2JjdWJuKfpXCWLCrxD9RujDLNTj8mhO0DV2CeJ2tf6cevBQU
JiFIfzEQ6WHZar0N64r5vh4O+c76X1kuRcg2O1sZbCd5EMmHe5EpUf6Nvl2j8H0nuaiia8WNCr5Q
ozTVNYmlFEy7HSXzDhPen+as3tEBlR5Z5DNcqnh4CMjdOYZwYKdlt2tMAfx0QMhw9P+tq3TJGuoD
CPm3AnVOfuod8VqM7zyWTyIt/GW+oghgSZejY9YUwYrZkJzG5DtQd2yzkA+2gZN3EUZZ6J/XP3zG
365bpt7Uc/UyVqHERJ3i19yj5Qf/ZktsfgXtNcpO3kEgwx2Nf5/keYfVn5TWVvmLhMhM6SSxjusa
xza0uJ/YpOhP1ksFcpjDpGbeMufbHDM4kX/uTlMX0YwQt1vXrYxv8rj/EuiilAZTBioFl/TBrqEj
0Uv97SWRQOGj4vDxNYYlxMPsW+5xnK4m3me+k6mJ+ZB0cE+ob6N/NVpouwQ7+xO1FgL+beKIwgSf
XevDLMNp86trQLD3VN9zFovWXUMS+nQ7y/KaVIvpqrg6VCp5pWZLYmaZ8YjSm9EFxM/w0wzq174E
I3N9DBp6UGHxt+gqTV1VhxqzOpHjXHoaQel+csBZx/bboAB6rkhJqli//g9cHGfxcGO+oyfgt8iF
HFcYBuwzDqxO9YclK0/UbitFcy+vbCp8ix4M0YDvjSbX0nKWaTaDIwLBHLLKBjEq2REA3O+Gpomc
WkV2BgQz9QaAKlhgxox9Rh/Oa5sjLYnxlbg9npKVn5LSlEJpSxCYyDAUm3sjEMCJVm/aOTVkJGO/
dXnapgKQHZdM991ETMPJuNU6CQNTIUeHH7oxY2TyfwGxXYrD+WAf/SEBi+CZKVffATyDvXRXInZ+
zpsQBsT7PPJIXE9uXtd6TK+BF8eRT62p14AR9KXlx+sjcogvPIAZUQTVfR8Vvp8NNuiQ8p865DiT
G8f/ucHAk3nntBVW7FTq/wgHot3VT0Ubj08qmMiCV5aRXOYwzWqMeQoWWoEcWxPmZRE1LCNwTcnv
O3+WzgMQGH/iBStg4B1POVr1g1agNiFlNriDvMrlDat5vrNAhESTEmIRdExfNnud3e2oYUafjbqL
daE5uccP896PalQqcqDUE1DBg2NbULexxCVchpwzVfb1O1YBCr82RY3ZXs7SKuAapPd8t6JCkG6u
yL9ETRBwtreQsu7nnjs9Lg2Y01s2CqJwBD6mXTFLbcWPPRB58QQOMukeOx6TF8tiL6afGdXjpiKa
LdUVxbmWGm8M8ESxwaA2enNsp1WRegf3AdZzJ26Mwop0cBNOQlGHeW/frKNmgJBqD20CnpKc+0Dk
0q0APxawtOEwiGVTPvfjCRDr8WzvFcDOv0z5Ln3KclOqluXqGZ+5bBZQ3gA56U+uBbtXOLOlaCzg
d2AkhrbWTLwoSbuxbvotSnQLVkrUMc0c3lJWVT3c20UUfPKsORPfXLAnDuBzJyXLL3Ju6V9TMglC
ZI1EBQNR5T3g7jlpN+fJKIj9xrGz81UGKPzWGdPzI7/kpudNkzoZihcKihUDzGZzo39Z6mFdYxtY
YFjKMh79V+lw+hNxQRTQb1Uz1ZpnwkeDQJ81S/OzXbESSSNs07LgAtBaklKqPyzdghaQ56wzPufH
I22SO7+vIVzRigilIkMNABBY1sJv6V+x7w+2Zxd8R47gECZRDuRb/18ePIw0N3hnXL0nwEELLks5
EFU0f0YkNLLwFuGu4w89+klt3tX8YFvpQpHldUDfAdgIgCqLX99XsvXZhox5v8ztx/ipA5+HKb68
WxZEA+X9cMYO8r7qm6Q14AnDj4eCtMq87P4jXGjVqCG832jNP+bsW2shjKV+vRmdASJVTMFxQFGZ
105BrI9RBjodAj9tNdkQ3Zq9zdTuClJcJTOL1m4JCu7Ua7hkKC1FmLHDKlF92LZOPMDDPoh6+cBv
wvR4/PCTm1LweduHqpu3oVhzupsxOurvZ84RhJABfcfaGT7h0ShR6ZKEwCLmVvIheV9ic0nx6kD1
9PTqCngGQT6iRScO+3iGqbTjJErKQ7vhdeJ/ejUp5/dWiapd818ey8Hjp0kS1nxCauL8+MFnbCH/
8IbwGYHHDix4Ih/oO9xvG0Db02DcGf30pj252TmZu9ALT66SLKacj5Mh7kJRI6m94rqSC3YgGrW3
5GQk+QV+h7R+I+iesWmZ9GziGk/xL3SXGYykjRl69qkZq35FCHbFlxIS3gq/x/OA/uULvyxhhvE/
y1F9X2gebC7lvxO6HddB1IwB3dXmJVFswppLc1oSgr0Fzojd+NtNUl2lGGCwQfg2JB98QX7Bd5p7
frVWzw5jfgAqwhoVtShbNwc3ShyvKUEypGNiVKbUUHhXP64NDhQpCZFdbcRDXGDUuebIe5O0pdHp
78x55T2LnFdiZv23BGr0US126vAe4x3YnMGDdTH3Hgg49X/Q33hhoThQE7fb3LWUOLBJF8NNrCIV
7d/Qkw5IkVULSGHKQvP7j/7uEwAvikDu6GF9hCIog6Hgoqc+m+l9z0o7o0iD2VbcDeaVZyfR9xn0
ATvRRGpzNzOdgJ4qyLfWk8tDlCNS2fe7kZmlynoToL2G2B4qeU5D++m82yukn35Cv8Vup0yKZE9a
NE88x5dTqFeKoy0kF5GNrfZZkWOoCTAWrvBfiNGcyGgWfGY8awyWsS0pGYpRFm4WFcBRZnsI4V20
gFi/M+/+fOG8ncw8miuQqVivNWi+Ol+Ua0WKlyEDLPZM3eGTqjNL2GSA4L3470hKRM2xoLl61kyI
a+/YyF2mmw6QfWNz9V/otZxzlHxoUAuaI758t85xoSq6LfFMLG2xhlyIZg5aK+O/4Sp9lVR1Z8Ap
g5p+2AfkEOY5v5OeaNHBa7hYk5fUon1gnw/7lC/0uAkB+MYD+ttQZdvaV9yOrJzEpONTxxzC+kvb
0D5ueGtVe4nFiJ5U7AYJGWwhDNJj41DIIT6X2FAhPIA/JUmP82lJKafnCviJuWsUlcMefmrv8Dd/
982OpgQ66lMox/ubXRcv+Y95UVxnCMDiDfcvu8EAdL+QtNoqnuzxNsaP/KkvrZi4vSPsrtkxOlxp
rftCmyYiqmJS1dfcYIuCJFP+IMOSV2yWAAk8IncBz0t2996DXp+ISwIM2d11G7L6EJ5Is1aLOMN7
cbYVWfjDOj5mXKsDjnheX7kbhNzeyLYYRdCkiCcUw2VMO/9N1QGOz1xIor2ydkwYw1QGc/FDETG0
q6WPVZnhgBhXbd86Zcwxl3+CxS3EMemiAO01rV4scM5NoxKKQKeouT3jqtVu1OteLLcHfTJlBpBz
vQI1LOZSwHet0QMUUqh24+oHEO0hx2WD6P9ZFyOmeHZ6ppYEUFymvtl7kkbzmZIovcQiGzqBaTPQ
H/nSyV2t1D4TQLEpB85KoMFPgpBk4/j9vojS5F8CkixxYwnX0O0Tig3T2nqCmZhuVQIRIrBkI2rw
truCyA+kkiVbzrxSwu4r+Lnxa11kNBUTKVzgjqIzBNcp76BkakC+DMLGoicA73ciiivBAOF11Ksy
W0lNmu7jlnktq1gZsGqXeXJYL+qa69ymzOHuwTl7R+0oHCScw4EBR/dOAHjyTyBXubGJB4XtrX8M
5v9qrtO1i5+wYJYmv9QxgrgleK8XLrkPYO1cg3JLzKJttYzIZ+GfmCFetYFI6tDJSz5FEL9xA4fp
kkeSoXUDjoZn1RXcY1PjY6SuW1ixHa0P0strNbJPFNbdd2YP2T6OxU3RPU4NK2W1TxWGM+asmdw2
8ZfRyu96e2gIiUS5bLPYIKLtKh4RawxSJtzmW1Uv26zXA7yjRcorv0vCNbYx+RhWMduwy2jISxfK
DFVvvJ9A2hn8A7vDTyaEgQ3wB/Ujk93Dv00RswBj2iwU1dmmI64/qCl8gSWejDbD64/DKs0+91U0
7cMzmcxKUCO3hSgbczuBZ8vpta4H95tGDEnirfM2hIxXCVFOvlO2blpyhjDKcD6iLlbaDVODCrYh
rMvDHJz5DoU3D1I1yutzamabf0oy9UuxjxkCmPbi5Y5C/numRiMFqdK5t6YbPSokH3h0Sfa6C6fM
6KwaKQeiIQf9OWs/s8zLGjWyY7HFAy/Q4Nswhq7by8pb6SW+UF8eiT7tL4UGXuIjdMHUciofK2/J
v0I9LgIWqaQZfP8o80lT7X8QShs7sJOuM7VCUBU41912sYlfwRs2Nk26Osd0z5sQrMqwd4KmjYdH
JQQP+P/ZU8imEbLyyWq9PN2KJkcQFU2WI8PI5+67FX7hsYVXeznUXAhNHNeXGwjxBDi7lphQxoh/
V2bVd2U/7si7fbqE1CvMXX6JfnTMagZiH4GdATthl0gwyqeiudgl8nPgknE+yiLH3Owwxlpvc5Jj
koxUdTcm6ARx/vl0+wl36cnX+xIHzAnfvakci2lf9ErYQoA/ZqDpBALv2EdhHbFx1vCqCBMH0wqp
2X9bVDscweFJz+ZE+Zzhb1uvzNmhFlNtgVgsR+5G0LjYYLxdZKf0qxVBpPr0EdEnYkbYo5Af/6Ju
3GIYbsMaSNFF2ssAPgUyBknjta+pMZeHdJId7zun/vUfLiU8bvaWDO97duggAX06L2WGK6R2FEj/
Z0Rmossgo50U8OizK9PuyStKpyuvapGxGnIddiguXPsvCfF8j/0FeUD82cJxwCfmKR4IaSsDcp0S
puNCvmG2ktujuc+a7WRe2UfcOzFqkJr6TSkeqZcP9zVQd7FBEcCh8FEMAxXVxD/m0JmcQfWCGflJ
/8mN+GGaJFngCXTska0OX86R1r34xZvx3y1a3crVxq+HjHkOtuLpykJe/Ipx5F6BrNaEeYWNGLjV
CpNtjMcRWZ9OeCHeqBTiCfpAAuLauwbrOWOFinzuCpktBW9q+qS/mY66msl1UtOutwFz3Md1netC
eQ+m0+VoUxkjDWQATQTFkDkj2zBXRmukf4BBDZ1Avvh7jnjg9Zw82h66X+lZnm22YTjCL3x9zCv6
96XGlCpht6tReoQVSIWhDFaX1xcxRR+qvKqBCBIbbvb1CWVVt39OrtGv69KeIdEDhOvwcIr2DFFM
di622dmXb0+WMA+ivHCI8/d0wi9x/szEeokcjcYwIxTspHMSKuKyVnEyHRHbafvl3fZ6Lbmrfbel
LRUazPDcUONnjm5ilHKSLy/t3LyfmD8XjIGP+eqcwGuy0UyZkl1B1/CuRQ2SRx7cjiFj4fXK9VAO
B2ra/61qm9q2YgXYI+lVvUr3+mWhH2iDa1IahwLeTp1y5HnsADEKj5efk8mgDd2pPvz+2T1GR/9X
JInexeaNrcgrEQa/wQyEvzwqKQvv+0VlyTLlJ5ootH2M5ODshjdY4//82b1BCUwU+kHj2j9GHkDs
HOB0fRrjxzAzt/5u5M2XipDxvkOo2NM2B8yhtcUFzHm7DAayFQvYk+B1q7mcYuw+o7uiR0afKxDF
pDgPViPXs3PMjp6klXQUmb+ryZxjCDNVGr7cku2eoFAl2qB3JlBgwwDwCFCNdHG4VEo1fSJ5+i9X
CoAYQTfIdnaTgIFy7XDnXRqDFJyXdVqFyNMi7kFtcxWVPA3wDNrofIxS1DFEzimxJzEgdxA+689q
MUVsMyY0F2F9MVwyp66NpSX/zzTGlcDeuC9yU8tPwQDNNj918/5nl3057xPBlbbGeFiJGLMIR6TW
S4tUHfCF3/VTjMdwhti590QiwaTFocNtkCzUjFzMiGG5fcj+LV30E50BvRRVRBOvCe4E/5g9wJgl
6Ifk6wNabz7h3bP8zPFPTSRf31EqC2a9XPn8GiL2Z9iTc45/DwUjSYxcxKNmN0aBE33n6rx5JVSv
5mgkaDi0JJW1IzsSYnvyyr5UPHa2qdYTUtPcnxv1WrnBxXUSfJyUlSYQbEhGbo5WpuIoZQvsNS2k
KJZ6mpWaHHvUchElKwf8I5EDVNDSCRaeh7bGVqCt/yO7JoY1th1NrU5PXDI3jluFEJIvkRi3sczf
CZ2ELfgdDdzJVaOMGY4Cl1pzEDdgsYesZeCVfT3gZmEVR9oSIJowQAJLjKaPB4g2rJZFQUnCh7i1
J0U1qZOWNANQRrTc+bym7CJGRhCby7SQM8PBFp8GAjS9xScX2RrUZtYClyqzG4CKUdh7Pi5bKPqI
8T+ERiUQHv7Vgrr5Oc7cudmX+t67Hkhajm3qO0ua6HcI5+3/9By32K/ncBj++H3vIrZLbtNZ85Wj
Ks69NWMBUTfZ4GiPCNFSTY5DL6FJWG8KxaMeZK4k6HLp3eeZkmL9Bxz89AuAdZ757muTXjs8E09g
yXoAS751B5f7KTU4kcUBT5zBI6Pbo455kZHhPquPvuBz2snt9TtEsV/Mmpf0frMxbJftC33g4OBG
GTSIdJ6ZuQ39QPdL2+bGn737YRZ3n1IVhkGm3kfvK/ZlmlSVOv8hc3xWPsPdf/SUp9pEAV3Xn37f
0VLgnojB/ionb4oYCZ9FIZQK0fVkvpHnd04lsbviOr3ayP1DagqjxRcMzn4gBn9dsP1JYXztV1tJ
AA0hwk87HhoT3jvGHk0d1so+z6ZGXiZaeacFcYkTKnhK0UvenUOplxB8Ei64GJl4gplAK+CvjN1C
Pxx5SI5ZD4vlCUC3JdGg+r5oXi/Jo2JYZWamGDgL8TqWRM86o/VynwSCpulmtKYjrCfi+Hjvf3V/
eKEfRPvtKPRyTwB/q3XEO+yVhlPCt3k/QtOUB/3hO1EdMsUhlcBpNOL/+t7omFhvSHkI8svbQo7P
t6qQjBmYiC/JJ1+DDmezUH3hmzFzBZhbQYiXRm866gFloRDPtswlINBPPsKktUX2oJDGvbk7V+Te
DALc/YiLbYP5Ss4O6eKLA8Hcw6lshtQg+3/AAeFwq4BrhDV8jKh+HaX4bLog2/puKs6HK+xVSgFU
r0DlLGPRN4Hj7bQ4Cg+LDbCKN65J6yUZcgmDWjtC2rMVQF5UepQFjt/x71y99emMdNvx98ADpVeQ
Bd2xjVuFBnAuyc8Nc/1mogukk5PZt+dwbGonILnbiE2mxfyjGI5TyHUaNBPND1HwDlx4L5HqhZmV
MXTt8G8Bvv2xqZ3lnaYPFQGm/a7IdfvbHKfZ9Qf/tRIeopapG7u+l5H03b1aAgloL7Ihz1zfHew3
yx2ksuXvAJq4+sPM28ATNGifoq+pAooJaer7rqJSyi7aEFXu/bBlexuDNiVgAq90CUAiFVgvAwmH
NljBq8RMODMaMzYFUAaOrFoghQY/0ZA5T9A5LLubs3UVZLq9LndL5JAUoj5kspmSgD7M45NmNs0z
ppvK2wkIdHSCle4alqQBATFdpZTlS1DqI+vWUm1m3Ln2U13k9lg0577y473e4PCEhLC2OF596Xr7
PXB8i2FE3SEiUP/lhyNdZyIGj03AqFxvscD3U448YC2Y9dplNFaIEw7N129nFt5/9lxvJN6bAk13
eWrsWNAwZVpQdhYU1gIcTTjgUGCzFAq7q3m3N/fFbxrp2JQE1XKddTZpfD5L97I81EB+Z+MyNXQZ
JwbkYKJ8bQ2nOGBKIQgFjLjm7vRUOxhq/Hn6KecPT28hBXzDHTtonqgowrVOcFQQ7UzdoWuL4mLU
5mOhI1VNX3ZLk31KkOtmodz/nMRqEq1lZTJ0mJmqf2QeotRr/dnkBBuX+ez3EFD2PttHpBM4UkR1
ebz7g6TsZA5AcjknMOj+9Ih2SfUc1tvPm9T/Obs2GqVo0hcAPZxM7U+8vfGxm+1aZGXDHnpgGXLj
WXuk7hNOTqZFYMRBezQgevmjh8AXLCD1CggY142SEgrDKIpBULEwLKR29bk4VgUIRqExWAeG6JlH
cBdgFk/1yX3CFnPxMBifeyxqTfHl8vTtfgOAbcMDRRMpKShg0nwOzKu7wu9OaYYXIE5Y8greHP1I
1vZCgF3HVzQ8nyANrKVhhd+qyFDov1/jpij/rvULBoCyJkaMpT3LzW4gwY+v6ZD9HBMtROYB53zc
KJeI06SWJllLs9RYXiMxNCgVYtXU3bn1t4gJbkn5n72cKXIFukAnWMpxhY1oxqnPd//xaSFsdUGw
odGRyLv9XDsumKNsK4U6RBqwMPw3gdS4ATwJ3IUkW/lKJno01pR5gf3unqnuouhbWaKd3zZawzwH
pUe1iJ95f1BVFZd/AtUIQ1+JM2l7/TPfcJCZoqd9INpoJoPjn/r/U5SMid6g7awLudifJqvjzsSD
XITTBH2ClniQDTdgv7J5QhiYpmOkq/T8cuoa03nW3Cljz55sX1GScV+edQHh0lXDJgJm69OYxrOl
33nL4x8/y4sQBf6GRWZoeklx8Wp4dckHOVDeI3p+xPwqP03lYKXVnDUrX/eJUpzj2q+RoT1atrdC
N8qJNZ771vbH14HoJv9ZuV3PefhYG8PHEk+E55vY1l9YPr5dZAhvH+FWfkVd3YXsiDbmfNIvAbe4
vlCGJ38fwOslSyWEnWMEit90nck/t5c3RslAUbLkDO/LuQzLwwSV9zGX8sSq4qSnZ7ScWwUGfmDq
Uzf+nzd52A4HmM43+chIMHhQZ7iUocNUY6LVXhCtP1kgyHlXPRz/Vjs5NVQQPFmKe9cmOFnqaq49
OBR4FJEnTNST2b0KSOeVyBV3hexeQHyI4MZeiNqT3b4CLKeQvUjKXDwZwdUQlfh3gFXbbsnmNKNv
0fqiKZWT/IcOBHzJU/tgS6U+r5koWWQrnsTLcXI69iAmpoVfHRz+STjnN6C/wbEcACl9yUbnn0Av
rb5mJpYaefUfuiScle8xUQgLXOtUmqNyQSYJR3EaIEJ3iQ7JbD927QrdIzGzr9Phi4HV15LC7sm2
Kcj+8Aq3hz9RJPH0J0jXplWhgo7gMn6mqpwIeSAkrqCNAWO3z4kTQMDYa9HpRUztVC00jxgt1biS
H4dnJEAHM+fYaS6KFpHaeI9RgOPVggwJz98tF5me1PrLpfHTMKOTblJBKqsMLS/Gq7yojIUx0IEB
9PqdHEa034GbahFcv4cdybQm+iAQHO1y0Qf/tI2QkdzcP70AhvHvZ1pWV15oxlSpqzoc/s8+5uLr
VUJ8Q+/ZMrU4bxtgPz2z0pCTTUX7t6N081xj97UHkNWfsWTA+8uT/EITNqUY/jHUkpdVOcwKfjrd
B+zD1DLD2j6vIHDe05IFx2EVJhNGIeqRymp3XWiQm+LJpR7WfUg2j8eUGir5MyALct1+ZtE0uirK
EKJ+vLEqhT29h7w8eKrJa8bt4Es+p891J/JXI0UgB0Ncj5ccdyoEcW6mvId0u463FUsZFmttRMkB
/NXiq8f3s1NVYge5f5UIixWabQQs+vorxOG7aLm5Cfmqj2Z6eoeSqXdmk5tCMD9sjY+Znyt09JTP
8CmU6BjsF9roGrs+GByFwP53qe+BcMsjPKmpqPsrs9AI2KvQdNskOI8+C+nm3tvTu3Re8vsjMT8S
wB2O0R8nfEizbbrV1vmh4k6tIteJrwve8k89Mr/Y7xQxVmN9crrZdgxjYGnXaQZ/tYzU6+HFoYyd
qjJaVqG3V3sxtIP9IyNPz2Rrk89YsCk6f0MejtyyJfp7yOadrQNZtfLilnJNISXzGa8jtiv/2Gdg
rrXJD/rdtbr2yrN5/0wOMWou2x9vpD6QrDiPut9fgqEtvKhE1HfeTuUCcWLm6XpSKT44FKBp9L52
AE1CRv7M5ORRsaizuoGN7OkBy08uO2NUhc8U0OArLBnRDGt1ev4NtrT7bKhbkAtuFKfPzkmfADvC
7IOLFej8X/gEQMfdlcOvMcBdg2oIO1l3TxsqJ/E/qfGN9BBrFa0ELzlDBT7KyYOek0Fi57VUDAj1
IN4CZvSGPBh2YyDH2PZAigdsSB/dIUrKwPMzHEKRB1+tVHdUGbHjqt/WCGZY43i+bxtdqOWRShOc
7/ZO3nPf2ZaGha/ISeMT6171gQaA6n3rV/DtXFFyFMe9ruJxhQBAvjhE2s+ATLc8uEUXUVmM+rKE
O7MtlHi/AszdYOxgkkewfrW7IhTE1JVh8jI2w938QD3OLpe6wFWzLnvs7aTnIQkGmXh+igsTC8tM
JkaDgc1LoIoHHYj6sAvjcOpE0GOQTsYBAQ7gBR8lqhg2QYCo1aXqVltytjqHJB3RL2DGn7LZsbo2
RoRcAAWWxhZO5wVBkEek2lVe9grNAmubeKWD44squ4vH21Js21rTttNvXfxckj5EIcZJMdLwwQun
ewBtXMuhbClMs7Y2rDkDukbczJGguhzC8DRBDPXhMiMvf2R8ykrJ9C4oiusAP5wUDdZrBEt/rUqE
/bi8q3MLblUrnjRtn6lhYIi9ea5E/ktr2p1PWSq+laqFNJDCVR4ukAkvCwfhkj+hXx1XWmxKrZwm
ODvUNZHlOYz8OLtfsCRIJIFmmglA4xnhrdXenMMCUZ4bU5FFjSURpk5bmbFwRhtuKvz8B9ApTooL
o1RM01cv8aFR4CWa85YuLGE2jrx8Eja0i3yOlnNyoHkklkorTKdXKbXnrOAohliJW2zckdfjl9a8
qLTnYU435DeYARhr740Zva4awvJ73G8yIGg3HJM8JcdZYnUA5bdcvrrtSEXtQAEBX7zjl6BMxdub
4pljVc7hqs2rHFuAnXAIw5dlWmFzXUzu6IKPXDUjum9sDHg2Wi5Pd2Fe8ygw2SVdNCpQq62hxOjA
7pFa+dkZWO1RuuInc2Dy9EZR2oCd1m8ITVo8OFtfJQsCS9K2Iedoh4+Cz6+HbinDVoLLSDvfYf35
r1APulR/DP+OKCFALchTbp4TKALr55f/6yUhVOhBCJIxL1CHfl2GkL+ejrFJO0yuqpheH16o2uoI
D2yN/0QMH4y2OABgHXMLKng3Qy0BJ5kinhuCRDwYVzh38yfdZjVSxYVsP0GpOOBGcf5/ZUlm0H8B
3b8DzaDQf+ESUhsCm37GkX6Ux6rd3GOFsTG+1tJ1MvPsc+I7cRlzMCMiHqOY5KMAUTRN6FVSsSM0
g7OcNovTb2G1QIVzVwfKCrSoTk775A2H20jIQn0uSV3eaoRPaonxqyUZ0gC/wduc2yKIuVlF1v+R
pragkLbFdXlkCnCGWxdHhpvyGsIwCTdTIDEckrR8bg03NNtueRYC6fLIuK1GvGcHTrKQyDcwl484
hg5BqM/XTL9tNxCnwnvYF4l/+sczYM+E0j7vPLy9EbMmjhXU3kpJ15SM1UZdNh6ZphhQ/fcx8oqN
NVZJHZfwk+U9rUjsS3bwqN8KWWYt1kq+smvqkvfyTZtufEccCDXA+euq9TBZlAQp4nku/WNuLqjk
ou8dNurflKe5LZPYH//uKCd45SHc/GwgjCPZT5k80ZO2xTXuEfCFgRoTA2/pmIJZHvN6h8QK2B/K
kHiTobKPVLUJRBww08c1v8iBFIhNl2XnX/3O3e+jSerJlPfEHVIoOfsSnT7n+/bhvMFCEinnTFOk
F/X5uCBeVVTlvIPnal/qI3Axz50ZOm70UB5xHGc4Vjx316rhKb9Y5R3pEc2xC7Q3AeWv8beF+e8Q
9t6ybx9m6R6QM4uQkzC7/Ylos/Gs3PE3ewM5k/Enr3BIVQ9qlKmfV2KIoHBf5OyCNPg/56PIeTOh
8hQKqIGzwA7ckrHPckyRf89WIDkRWV3RkRlcWxzUGqLPZPmdM4e/h0VGlSfrPEcm9IbAaGm7S84+
8RyeKTcACfXo0+v3OU/JUmbNipKwIUlSyG3Yh1xzkWwK1z+MbPYrc75V7npgamBXvbRG1eubFilR
QwilLegMXLgr2FIYK9bR0vWIWeJkvLqaVd3NbwYonIiugTTxREZcSY51dvsMTFwVyG5Y38FKOBeX
bcxvejPt8EzN67IUrRmjmJpWPF9Tndymn7cLccL5dkRyG5sBqacsJFdvHHHlFrJvKVnjKiJ3yKnA
p3CNhqxzuXnBEpEL6BfQwF9IXDPHorI4Dg+airaDhyziyvUjvggGaV2RFeYnNu91Z9pXCT97OFQj
jRcsPJM2jVMhRg1NIqV/wh/VuE694wHoxbcIWt4gDgvDLrNyrlJKfGmJm0SwDyLjtqvPCrJs5rJt
hw0trTOhcGyaK87Moj2kRQ/5JP1tWSVVDhTZWZoufycV70DU+owLKWwzkeZ9bhJBpGjCy6I1xQcs
BKIfP+n3yiV4jyIDf2pRqjsCbc+D9zyQghBsWNUe2L+EP94P6VKrWC8Tsy4coffWYnBsxpnJa34F
gqel3n73bF54exOS+UPTc8vJJ5WiUO+Q+3245w2baS4T9Fga+2WUo9SoJdoh5evNDMZqGhsdfFNs
nKnTLYc9pmllG+a43P3YpogHgaBO99OOhvp+4MIK09uSvAnvf37jl0oXkpQpcmVTbMuA9E2ml1iH
GM4DDjZgzsktt39ddDw/dpLL5JNhz5DRpf0OpsmophTOSXqm6HMQdJl74H/3XvX1viM5i6U/rGjC
vMnaSFzjYj6gqBcsNlM1hL82IVu1jo1UYQmJe2IvNbN13ujHAmex9p05ZULp7SE06YTnrgccJ10R
hLaXOC9roAoeLM7RYhzEiapkt5SUyg/CH4Iq7K0avOnHXuWX8k5fkqHlRsfGQJrqJZsaPQmoyFj9
KUWeu5cnKFGUJGNe3drT9FQxi7obn8g/hmfu4gw4b8kKB1ChExTgR87G08WoQcvnmcv9z+V0XoGE
+YMs+zE5rQYe/jv1SsNmvnN3+oiI8yH2PckuDN5+paEH2/cMBjurI6RGwAySA8EJZRkMO8JUvrzm
LFliChjud0Tw/Rw1hZIdR9d1nRiEn8mriOrHIC6dVaSIWJzh7U7D8VN+fXohNufnTEAig9+xJ3/u
1dISvfopm4pxcxJQe1gdTj/TYSC+erRf1ldHVgt153TvjYktcbS2RiGBz18yJgdNosq/dGU59T4Q
awWX3ROwSFmngqM/QEqAwlaX9hIxlutfYwgbpa0/M/k1hlAx84EL4vXnLBaDCxF7phdkRcDoHSAs
whrneOo1L9Kvkv4WudclHoe2XYdPZeF85ZX7zf8v51Zhazbapqa1BdeGNBDgmOTJ4wP14I0Sy93x
TXzq+n8wO/ni9SfZWRg2gTDaRC5ATFvSoYi89AvOHuKPLKIMbzFml69JOAH8xoysj5cijwN6KDcI
YSQmVVsOGGWtctZd8ePMcWdLDy7G9pSTsIR0nR67FGQFegtf2Zl+U8HOKhkvvtodU+uzWL3Appwa
vbgaPIlsczsUqesBHvr92Ghml8t50Zv4qpdj1psvShAHoaW5qJpR4N6VMwT/kF7EBikcibTdyc3I
LdVvDpPWK1MpSCMQyEdl61f5F1oo86GOjCP3IkbK0u04k5bnV4CeopBGDCa9l5Vce2sTsjaqM7l8
uhKsVGhhmj7XhoHnuIy54AYRVTqJeV6oQ2dTmLESvrumoMwY+B+PKy+656muHEA0KLuoPYjUKrXp
MHNyWYdYnpiPtB80LMRutqMllH4CVmhn6Exe8oE1IGdFwK6UeTW7ortYxTAO9mRZpMT0hF2PMAYc
cC1WooaPTOy+zDBrt2Z0S86gyz3YjM4Ig5TkrgpSzxb65l4GpLBOQxPZyVPC/2ZIIsBYC/puPEIZ
3ay2Ez4ck9xNk8fCLyg6PQTDpNBROebkzlUu+iYIIJwaxHvwR6OlrdHmnuOOrsphHcKQAkXrP7iB
ry8qdvi/LnVj89SQ6xEGGK/8uuk+NXOQ/ivF8wA18fXMwo2tcCUP/E0X5JCrAl/JIxKD3A/wfx2D
2BNZ9dSe5FWqdkcKeXdowPKemzb8Cs5SAXj1hVUOZXnOzViscj52wOr1SLtgtuV4lbLW7ElTXAMR
+OiIx3so7qeP9TU3ZC9D5eK3ivSTz9lCbPXZVHlf49AAHdaat6heffM2/cxyjSAegBjz8O/B+ngx
Au5JyIT1ffE8bB27FzqcMc+4XxdOpxoF7gFx3FUG3A4yC/gzkjvUllhlcskyjPcKNnNT3OWUP5py
2dAzz/KYsrllYeBn/4grmmqFgP8XFadwU9mo7muDnkuGNzQip/2MOFZrWpB0F6mv4auT0sydSx6y
aprp5hnKHOjUdlyk/wM9BGK5ESqMCiFPkqRq7e7KFjjWJap8MvBUdlQEHokW+mOh1hvrTSOhTCk/
VN77+LWOJqEoUMKiRvFZDSXhWnHd13Ss3UOd3tfTbW39xLMK64NZ1JrIiPGfgUE5nLhcPH/Wp5XX
hX79bmVAc8f90/Q3rJRYd7rUrEmyvLgJR3pJs9qt7EFMyiafkPxX59s0vNaeIDU1baYIzuXBfwXG
mGybZZKlhe+2JEPYEVFHQFD9FzxF3tWooT7KlNgzitQn924IznwLnJKCHlxJsR5nIWwkeMCsEg8E
EGZS1jBUEcfhNb3x/KiBngq3sq/4oiydKyS9UgWFlDy3QquNHfWPDuoFd8hScgFnmWickce/qp5I
cPJj7QquCDPoRMs6buoQHWSjq7qUzwqjwngzdgW+ai7fgjrf8Af+IXCM8M+coIK8RyuO39ANXI53
PULQQp8+uPNLPHF7q4o9FK2TKefQASsbUQOLRZGWgGI0wQUw69xO7iYlxoI6huTtE2bPBAx8vNeJ
M8o6TRX/D5jeIJCZKRIeI7RCGQgnPs/53bMHcX6juv6y2cCXd6FE76tyclVLQ7f1ghU7ix/zrDqx
SZ7jUbokTazcJVlgIjWl+uleLKoKWIa73sQJ3Sh6JmFk5ALyfxllhnj4RtVGBJe46vH7nrFUqb4Y
WjwvlPR+rB7pYeAx6K29tqt5twoHmf9gQ4GQCv+SC6LL+8KP6yPdu/eT9GmAEAhSIALcSQeKchxh
+cvkauIjSo6K6Oxq876Z9jBCnmrS4jl71lL4vh3YyXVqTdEuw8B8M2EqJ4ggR2fiAIwlV4HKjcW+
x69OGV9hAteKKL/s23VZXX7019gYerVWstb6/IoWK+C1h67iwCtcDUBVlb4HX3naw+4uBQioTpgm
8IOoIWiY3cqGHo0daypCS3GyPgOHSOit33BA+TKNvjZAszaxckbNlEiaj3zcKnFlPDa0k7dYD9UF
GV2o1VEq1e4l2kRLJmHEIU+ZkNxTxIZjcNWVhQFaWZG69hT0xH4ZW9PDj5kMN21rHis0vvwxyKhw
Psm2j2rIkJPwexvWoj9B0rNiPz56Z2HI8y0o+C3ArEIJOwRAlQJUjN8t7vFGZxjq6tKgedrrjP4O
MniAKGjp2grA5n6NHqbqAfYtR45rRcS1D36Wdj2WcJONatoO2QZpAY0dUGzjKQpZ9WbNp8qqUd8p
d5PFzzd0TNTJrjaEnfm/MR9fpv48mvqwdMgHrPDBOyIThGscTAJF1dGj6TVpCaFdHVAKuLOFEUg+
ZJNhJgbeGS7iKLunv059gH72GulaRFpSoaJwH56FHsTKBV+jFGIoR/AMoB417S/znohxlIFno7ha
/dxerz/D9iP7jEVz+MMO0VI07uWUt0uVEpd9QkRSYxyN1IUDc0c8gMbpYNEB8gsFyPcJQ+etKdLJ
j4zd4mLWODwMmpQoRsq2aG5VZ05xDl1+Ri3q0kOCGKtyJJlbZ1hTzu/nscyJLCKXUngs7t47KeL5
FE3NatkBgGeuH2HdWw92KYf8+dGXT8jZN3gFIPoIdUWELtIwKONjZBBEYbWLKEE+pbCK1CXMjO+f
YEqWTIvS4+uQK2vwzmZkyCefM7BX4RgRCPAcGssHWbLLLzc5Xuw4P2BvYVcHuekpuomzNKvnlfUZ
x/jtIKTzlyWwIk3CElNAMD5I0ToFdVxm/Uh0XXO4UG31K36k032tDWGxxALxAQ4DfuOj01vy6MsW
5l8mWta5BlvFXMwXfKOq105Wp8Wpi8kuCKq88PnQ5I0A4Q4Ym9dyLQL6YJ/cDCmmVu+rCtCwhO0G
tDM7LUvrpYEUgnGO2QC5VE3IZu2YzcZBFK1YGbNXPbNg90bReFXkPJEwynsGBZ9NQovLJJ3Jfauy
eZA/sJz/DcEP7OzyGW369RbrHIpF1Uxh001uGbRdPj6SYB5IZf0Y/3xjepglQ/SEJcaohKAn1jG9
/CvEDO1q/PgC/IGJY8PAmCh7xwp74yreDzZa4xlbTuwhF6+V0XM7VWKXRzp7m6x4l1jTicJpUvUN
SAEgwKCdO5YGeOGaNfrNHl3UDNH6mtw/kfiIqMRM3FMc76Q+RNXDYMzsROKt8gRyn9cky4K+4LBo
0qltm3hlYDO3QEzplFOR/pQRS+nc0CqqwLdWc37WeX6YOLRqr8gcG41MC4Mn6xYycfYr1d/v4NKw
Xomg4Cniji0dwuNo6Ie0newV7amkWXAZXsFRs/02lZmeqvJjgoqMNggLXMNrNyiocrsdGQ01mfrC
ml98hfIZDMmkz9giIU7PRffCeEKt9NTm0ECe+8jgdb1UGob7jDBfvC2KcDZPkHXg7PDJ7yZx+I37
Dkti1aixRNUIBKvhQo00twQC6C0maf/hPrM4NpWjki00G9FvC1FPuWILZzZ1MGo4hpQQXUIxxeGK
OuOlCdtmQiMEXOl0l7kS9Z7q/TLOb6+TCGytIIn+zq2L66WSd9/kQh0Ylgposd0hGSgfED3Z69tM
Dffon4AyQuziAx7zChBIVmU5K4uPk2BKdR/YlQIU+2rLc/4Xy2CFYxC3Nn5WB4515o4DM4Fec7Rf
jjiRjtQpwXSaIEO4w4GGS3/xKmhszYjeH/CdAYx+NOlCxP9ouGyXrsUHbweaMcfAkYUAh7kxiuoA
RjWJziafpgcwxQB76rGKRutADK+8gQJwQdGt5mxFXEsplgdd9OaTBDJwgDTpLVQTwf2Qnt884w5E
pHswtdAfAd1Zd1SbVK43HWUzrb5oD7BPF2sLqJ3FhWW8nQC46Dy+j8DQL+fivcdWKgGBMHod4W0l
8PuoBeaUs/PXf+CgnzWbAaxIJr3LiMuC+yLXx1YosaRrfMBG/slfohupO5Yc7/2ElBhi+0PHYbPL
t5VbFDRsLl3gE2ruTe9LCCKPQAVjCMnCwGfazsDS9HUqJARnNBz+L7l6MuxGyl4TH4uB1qWpZalj
UG0d2tbPn0TXyzdGW+YPphF51P9JcN0VjfiNoJv8ZY+cUiHOX7bqJ3PdxwNiOjQg+g6vaQa5ZYXX
KkiJhs/UAVoTcuULHG1BBfOi/U445ADyLjhQrgUkKQ9zrrbSuRNP9NbRdiyZCYCrCQJIncF/MaDv
Tn5o2pQiV7pm0RLWuDBGTuq7lGcDYb2XEQqLPveV4Biw18YKEtpinjNJyVL0/MQQ4OE4xwSmKAkq
4W4oJcVRIp9hjHoeQOcCkzedze9WF1qyDd26c+OD9dz5Y8MnH1owUaUFJGOkmyW2LZK1Mxz3iLm1
LcT/d1kU3DuIkFp5uxGWpyM4Kc8erJDzSLf9MouoZGeQ3WmyrpgSkKuZE59QY91RT1CaPlXBSAJ3
VLCOTCHXEeouENEs6R/+jVOXg7hVSxAlIWHeZAVMxFuZXlIXcvowxB0ixxsJ3JYmvWUAptIj7IWQ
smmtE9u+JWsTd72nnt3XQY09KdjbdJj3Xt0qYzMBqCIQGskg310FA9awx0yl0HnxU7FMDHnVT3/k
8CLgbskvZG2YvgIYHT/3YpeVyKUP9ZOQMLJo7z0Qe8k6a3Ge6M5IOxPSP/2IWkexFNgvN0z9eDBB
SKKeIBlI6MB7DOIdtNbqfvnxsQWxC9HqUnOjhngoUwZrt0/ulPuAY4th8+wlDXsIX7elEnb2Q4yR
/iAzRuPknUqg0ZGWA+yIUEnHIMr5y+A6ieZsNS7ehFc8bcFyceGJ56kgr/bypgeGyGtX7Cpljdpb
/bS5m3bN25KK4I+U0gMZNzpvp38GmdxrU0Pp3DCBc25De8n/MNijBM/mR8UgiC5Yrv6MhKkKRPHO
liN4ojG4y0gFRWOGTH+wc3XRFx2XrYf6k8tdM8MpZ6KlWWIZY0KI3Xjt1VjUaRmUeGs2mxhZCFiH
jgEAktSKBGpBTltsDeX2Yp4Cccvt1NF3YRtTjLC8Fu2WHyldTNIxFabVwbGXLlm+6oQ3rZV5PC9W
WXM8XRso63lGxCzDjvV3wZr+ztzwjX7Q2YN5FE8XRySWu01BfcA/Rq4TayaL2IwiX/3QZMhTkd3F
QXBZgFGG7PRCFFxdBPnJBkw+OBUioLtS6fxz7hAk/qcH0ZLxA8UUxKa5JEsQJrgJfWPFeWfDFORz
9oB4PXxJTYfbcefZ57rssKlCl6TSNWaf8r9eSLGsCXEG6W23Y40d0Ne7OZqnkmjQZ9rgqBxSqq0b
ypObPoHSGemGbpX5O770ZnhDNw98uaIYKv6iUfsPFAT153iIGH8LlU177n+HqN25bTLLmQ/zMkEG
SwY/yCnbWgHceGMoK2JSmh/5QWCEO2pVrLThDP3zVWan0ObBOGaLWOt4u5p6CbNnyTPF8YnFvpNd
0Nf15Jiq4NSlt7TepWYPtv0PQkPvoCj5TH/135lRjx0j0xzSzEB4RGAhCckbIqzFOuOP96ve81cf
AQeL8ldsK1pEXeQQuGKypMCTMu+4IWI3ljfMxuo2ogQo8r4YCcJpT6puxrTajo1tjLDsnQ5lwLuy
ofwb4FGQsmMS8KoOtNvk0Vmm6AuS3Jz9gCiWy7RqPWWbbLA2E51ehEENMhgJyO9foV9Ded18Z3u9
cwZOwvj+ojYlmUIQ0gRpEpVZa0ryRolp5tG7663gmAKRpJz+ghv6yM8dwXBoVF4/s28mPn0dRTCo
LHeZas0440WwFTciAceZ2BL3E8yRrWOu9dAqfshCW0JIH8PlXYs/Pq+FL5PUA4RAbGd8D7XUuJMb
5eBZmIAx+Gah0BZgQy4IZdRbP+bpzcw9rT7qgaRszlYNQ9F0z+n3xdQWO2I2icZlXCZ99XiHXzUo
Q5QYcmkjYc7JFLLaVmqyIpf7fc5gWWVntORCB86SuGeEdJ1re1T9qJXXB9QkVvG+2sctILvQ0B2W
h4PVeIBR0TnI+e1g15jMpQuVHB4+rIF6dYi+1EfgEls1anC3VyYENZY2lVN8IDchkwj6BDWE2EAX
fjRzlydCH7QLAufbFCEG+YEW0pAknH0OyQthg6tS/wChJHShHALl7QEei7zaADhpQJIc71SbBVK1
8/K8cWniS2SjN20znFLRBp8ydl/AQBWWgS6E4GD3/51ONHSx0P+sDkWjMyVZDzbMQqrf8iGhhp17
uc4nvHYCMCZcf3As+pyhgI4pg0hGjlRdaTAcZf/n0+8cyj2NrKy2hGvmbG239l+UX+0Z+T9l9NnY
hW9iuxDJR9mmsXtorueE2OgSazUf3yI4wmyySdeKBa9bUpjEikxtiXowALcX+qUwPK89u3DHF71i
pJ+0UeMSz7Wb4zUryCxa75Ytzc7vGJ5+Kb667t3ontk/5X4dk79heO75aFPc9o31WDckzIwojO7F
n/T6brH0SCUZWt7Ke9CDC17htwoOPbvlJVILqgKs46mTkvBsQTLZf1kENp3fD+jGIKCr/UVo/E4N
xXVOKPumi1tqD0J9CIO5OiRfD/G2NEfh1mMVBovlAgBOUiDMYQN5aor3CyEtQxZ+L0mfGQlmFDJo
6uo9cVAs5p4BNHWVnSwMzO18cg0hEe444K784Ej4AfKHHgdpFOZ5ZGpY0929oHxCRmFfi8W5hmxZ
M4yULKa5kGCg+fTv5vKnBll5x0Uv/v+npy3ifrowNcmzbXcIuNb97zF7rOsh7bK88QSppGTlztoe
frz+W7lOI0dqoqOunNfbmaY/6SXVnt3mUPnBl4CMRuEeCtXpVSg7BIicrBUxynh4oJ4j/hPDcZBc
gjFZSEyNfSCMrCshHWdgUYm/QnpK/a86nqjwyQxabaV4iev/4erHQBekjO5PHcv9Iw8Q6rOTF3tC
I2Go7TNBdqEd9LHfDtvQGO1KYd0gucI5YImHvAEf3B/IjmT6UcdUOv9SFI2V94aqVal0/BDapx3d
fcfRCo61I4hYBtQ9SmjmaPHwuUfv+5P+4D9O/D54/mH5Ysv97HVxG7aRdIjHfZfv3soor8059loF
iZp9gwoNdVHLuH61TEY0kchkK7VxxPB5ERL3EnGZ518Rd+Yr4MxI6oERZOaP7sFsqR/W3p6A9bWa
JUKkcu7t+kn/mUB0cM5LLis5ZTahaPUwRRRwcOTYwyJI7LdRqKdqOO4ODH+d6XfDBOSNSDQ1LCOE
krPHn0Ec6HyTaRg+jKPrCnJjMu16jbDNHurFEmMRHNWXC4htOzGDxdhnLCgDGDD9kkfjp+dRsWqG
zBwbK2DhD4S4dMPr3Z8D+P9qAsfTQf/z79z0bV08B6v/9Gv0VIJMJyJyU6+TtdyxxHJ/UcXSHJic
3lUq5Am8XvWAHkVpfRk3dAfCqt+9C82Vw1ZLzaYi2on+albXU5O8UXOKEvJ/bxdHfc6IBcepmXr8
iLnsZ9VrEDT/5qy44i/Rj+khfWgW3y+fJAOZ7DiMMt+ez7QBKr2KyOOcaK/Rs7p0fAA8coDkkEgz
pSim5Xy3kykAO0/CPJb/gL0lzi6CavWIUjUhjAp9rtKZE8DPYEdqgBUGj1TEIJGYYQUqxpr/1HMt
PJeT62DgNuvaFHY67MyF4e9HlT2VVYp37ijB1YEZPk4BIpU/V7WDyERdUsQWtsH0foK8Hy0NX4cz
1anvj0htJa2c6eXbh5TnOjdcqOSbvMmu2Gw9RkCuIVELqREuXDSEx3LmRevWwEdtVJ3rlvBNSASY
4qNxHOJt6tUbGuZX3McO87JIPXjeQVeYx5ssBDpktxAB3AqVGcdXfKBu3hfHmk0sf/MaasYjj/Kl
QT2oXS6D/E/Uy8bhTEI43DMxbb9tBYkPF3Q9H/g4S4xZEcw9A+PGW04nvPAq3um0N2kbJLsdb9Xq
GdbdcJH0zUzlywB2ArwwAbTE6zNbGFn0RgeiiocSgBycFion9DhMkJuPeG6rWGsPdyZhkTPVn647
2CO3NRcmZQyl98v5xXl8/bhJ3gzltwOGMtCnQX4nvo5jrsXaeDWdimkuGvylftNczEv0DqaLBJ/K
mQmRQIdb+jn763cLJkk9Q0GYKlcRq1r5JEoxfApgYVvFERVoODvXww16rgkeAX39WF0GukMyVgla
TA5d3z/Ie9HLEoxQqodBcDUQApzFdYRwVHOGPDvgqVHGaMjJJhItqIhNT/QwMJuFleLIbC7VxFwL
kgw15sj8chk29pnMMjkCjFTyEVbGDyQhjWhpc58PwqQ2mucl8xU9XeeuEOdAAvJepNrRpRDSowoC
32wRVBfZ9ryl6zbDkiOpZby5r9wzXYgBkjYJLITcAoe1vSpKU/i2WNYrzlms5GfynsdCBj2M1Lq0
nxuevmSDJsbdbxKYIZmqNazswbRQm+22/w6V47pimXFKBEVLqiy9ml36ZaFp2KIeKFqIBmenJ2Tz
W6Guv5bT4HbFjRHlQE6e9ol9AHCU+qOt89SzjRZdcrd7JHYM1jzK7NDXK+OGAUUwD8vg/i7C1UYH
disFOA7VijNtnJy/FsLGjmZQaSQR1rSa21KsaEFIJObsy5FaYfUHtXtaVLQgrMK6/DOjbW1jJB8k
y0XZceyGEcZrpEJvsKGW9GmDBDq9DtTeiN0SRBBTpBodznF9nfO2EBW//3HwzCIObLnXzvPDCWNI
+bFaqiu0+mY1WP3Pt4f73IE/q4LTHrygRwjYPbrFdtuVhWKHFbgoFc6k8+3xU4E2CRqY+LtkvhxB
bPIXiot46rpRMORYQ3X6uqcu8jlf9fwe3cJTceOYy4QHYoOVFvY/PcsuC0KYQ1hG1rpYb3r0LFRG
i1Sxb+yo+9wjAkQahV0tdVyXCfvOmgDYt62t9IXnXWs83ONVCVEp3UBOPOj1vN0/wkELkkZ3KQ2m
FdsXXuSksQ1jC1PiWApxaA407qT4OE+cImil9QzUxxNbnRKpehgOGyA541ABAU1A6LDx/uyRv96H
+qrzVkzQaswJJ5OIQL+m0oPekUOpgM/8q5E68pn4uciB64dFlDlSz7MS8zCUsMfN1B1FjQhbJcMD
7v5Wn24YCOtJU7c8YCIYN6kVYJAmjOmZzV5ppEHUG3ljhvCKSS92X4huJTanoi7mHvWZG2PKU1l7
c/8TRP077WYGMxNb4G3jeUmWkjYJVvEqj8VBhEJ5NuTSvqp1aEcCWPQuPev6URP38y6gdJyTgBeX
fd+UIRF/motxmTzbu4mpCN4yEiYK2NEWVDI6UtxZx5i/mmqY/Dd5Vlfwi/nEUnwkYClMLdzhIu4z
v7SwJl+wvOtD1a660jnJb6j+58rdQS/t+agr8B2pjlACSms/UvXTvuPo0Hbk3qHSmKjepjysx161
87DpctdVJPQPAaSjh6+7ydBu1CSk1Ujo55+Ptr52S4f+yERCpY0e8BUhcHFnxRlNC0SAXGV5P0cP
0AH5c3ujuqFxw9brYlld0uBuUID5sj1ggxYDCRYMRiMJQahYA2f3XXnigIiiurE7RHoV8Un6Tdnm
RbI9Xfm6CvLVXhidZRCQGFrBjRelFNVYxE3dHMLm1f/YWU7i009hQge5hBxiWbM7otDPK51ZRwQd
UxgLFwgblQvF3wYCfrpf60Do+04NMKqqg34B3nZNZn9fb6vQ1mjo1O/joEnCddQkfTUCtrdjI3os
y8bC47Gwb7HL95NYoUucancXgQLZV9M7y46Wvp+fot+RbWoTq9wRSLIqz9AwDDqxW5YImmvYG04I
0oc71L2R2ySNtsh6YRe6FBaLUHbqI8RZ/nRQH6rhkPvHXqMX7iXDcfA5Wq0GYu3UtFAjcgbGrc5j
CfbpDnYzn5KkG3GgKSVwrzfgfui6q1drEY6qN5DPVet/dlTn9eVdBj+VxVOb0hJuDEr3HuzcCt3T
U99vstkr3Jf0juPZSCgKBX/08GySPx6eW78sxbst13eLmX5IGr9dA5KhTJfmT+8Gv0C5lOtd4q3d
sPYVWncWHB9ikHk8wgvRvjPTe/biyoXr36UqahCBQSXo0sK++5QxB+nJUTLGVhaiP5fGFNOWir1S
BQ5vl2td5LMLvcs/oyMOfuSGfwOKALHv1IjE592iBdH7C2WC+Bi1+7iZQAmywbJ5pZOR0fPVflnn
AJJOfSUkBXFJDtDXnCYVfjs89DNHwQfIAzawzGVngrD+3W1tz3TmMhnF/MjLkrw8YeQgGOQ2Tklf
gbUwupWbwLWsNiae14SvpqrHZOIWxgq1QSignhXvLoEQypqmQTGruiFNX86vk54cndqyDJrjL1LB
yS69uAqMfwsagx/wgOPy3uZfp9qIPDi278t+VSrRljcMZ8qlNAuiirhMafOG5qCBKrmdynmsj2jt
mHKdx45Yd5KrqyE1daE9UM7NDc9QJxlzYyjytqJmePU7lDRKiTz89+/moSX8Id9kNcK62Q8EAVaN
yWhTc/kCyzQg8+opKju9DrXYcoKmlu5Yu6ppqmjpwV9beCTM3xuHd4Pphe+ebWQZ1C0eDGt+QMQz
+ojOkO/ICEUcPZFb7flSbPg+IE01Zk/xh0BWB/wGqWH9cii8C2tdLSLIx2xEswmJkdv1xMZqHzLq
fu+3JB/LZhPDBVsqm0J0Ia/VDc98YDgfUdxw3KJszxAgM6P5pu3feI8r5mGhI9CiKPkHAiSVdYiu
eWmBo4v5+epRqNsIxLQ9Zas9SmerxYBcas/BugFRfBjaowpqinVRcNziDecEL/c0r8Fe8ThY4ecl
wcou+MWzFAhNSSoYGqOC/Yh6ZnNWzdEKU0kHbkB+sC24XYlt1/SmSDTUtgVaaaWlDoSPpqXpVyT1
Qy6Ni2VpVaadArYYJgfwgmkuLNPMBphcbB/2lE48eaMi6Qpt5IH/oOjFSmSiUOXXhyldK4LPyxxr
Tf0hH/WjnWjy2bt7If3U0G4Tu9yEVGQLspsdjRNSHe2loMjwA7IjLFls3wZiqlqVA9A0rpcNljEr
SbCV/d8d5tXLhhkL3TV4B/ZioPSlce2c4vv+nH6trFDwA4TNXhJbylNLXpoP2vQEK79G1CSE80Pr
CxGQ5r4FsFJzwbvSxLonNDNWU1Vi4rvqLRV+QDrShAcUheGYk3efElbOiBOaPW6C2mE0WOp91Kig
CMipIBlWYlo7p7flcGao56NFagCtr3CgfQkpUHUUPJvRlNEg7C2vqUTTYmgGJa0ToOBCWf9oFh0p
qYulE72V/pBXL+RLbIXrf9JwJzpcDQpyL9IToN2kEKbt8GObULU7o9WLKk1lIfwycxkzanmZghvr
D28xQFMKaTR3NZPQEfZI4QKD6JNs6OHtT274mkE39Etc8mjY2EsiZ2cnZZVb3inSbwFkp7VbRIsZ
+YRVaWHtpZ6nfh7r2W5xLeAJJysTiMo7ziq24T3rJMlJgrgbQ4haLU+HV3qlKzDn/ganAEBmFCqc
YTGUqWYjgaZ6wjIon4DGiedcQuq9PmLfKFUBt0D5bB4aILf10gMbUVlDC4YpixK5u+NPTTjlIdOJ
JseVvUenw5DaQ6fzYbspUnbQDntg5Em8FRdZ4BVKds6+cT8Xt9s2lxr5c0JgLqrKAX7rbtFzH1yx
V1se7oru5No48fFkVyD590eenxH67aHkD8nKL0SZxFEVIHwn7oQ/p+0bmhmpox2Mvk6rl4J7LBj2
9x75sCssEZkw29Rm3lEX3gocSqWQWomlSizSNmIByrJBVM1k0pog4RDl+P2EMppcLuGzG7lEtNyU
Cg1FWw8SEA3ATVqbSaNhHU60/X1jnNf7YwXxg3wWw/GIzHR9Z2LxEAw4w85Lo26XBr3TJSqqF6AC
oI6VHnhlzQUh2KQkrtQ5u2kWY3pMhorNjd6/mEWHh/GZQaamztw42w6jHoMHeM5cumBjj36Tc8A4
ZoZ91grlAzN2AIRj/7BE3iyo/zlBRG3tFjFa4ak9c7W67SWDiJiBIxayNrfug30T6byKIpTzURdC
0MvxGjVB1zr9GlH2n25Ju4RhE4B9TttykXg0KzEKh+1xF9CKToRR1LYYnYm+l4FYX2xxhCZ8vr6z
iD7S37Gu0dHv5qc6x7CCYW3pe5uWhntKGBVy3cNq7R8cQL2aNeQPtdyAm7z2JKZrWbMhV3p7VYtX
APTw0QHafJ0Y4dsXEYSDWzz9T5ncpXlgnraFYpE3YBYbWZIKrmHJpnb27MbI+t2pFhqA94pDcxUm
Vc9aw1QO4DsnAOu1WnxoO5feshcj8KUsmcguwrRaxEEKVrudoj/XqAyprBw0CKB3EcP/JmXli7Kn
G5reRmWlQaOAEUuiu2zTV8TETV6UkrJLZRrQrtYNyrUGp9p9bU+e8qTCCkqXklDoSWg3Hy8q1ppR
A4KaXZ+11kZ+BPB4aR/dlQdtptwD+KLvPjdRqPk9NB+U5A7I88byPwyCPJHRVbjGtQCRsMl2SbD8
fVAnVsNBojVfLCiLagT19jeZ5mlgoPZuiYi0JK0UsaGBBfCrti3rMjOfaIfyRWz1Ac1mGypLr3tB
Ryj1t0JjLdvRTuer8iM8vl+GrDBv5Q2OI0MsCaFePBiRYJOCr4I4XL/9wHFf/qu4SmITACEpwmfq
pdW8zRrtqMqXtS0KXPaKn+fYum3de0i+Rm0hrDh5gT89tf1YZxui5UyD4zivaRxjNsLO0e5Bq9US
TW07XxHTiMKDfHf7zijkfL84FCXWkpxxUa/xIuuNzSq7cOcIQLs8SYvy6xl2bWh8niIwjavMMP5W
1oMQGrhaHBjulR8/rgWJ8SV/TAiunZKCOYSue2SIPujQW9EBE+7W1tWax6u9DEns0f62Im13Bxd/
eYisvbS9sPrWyGv90/U0R0m3z4hL4a0TOBSVcQXhNyrmndX/wI380DcpDbIY1o4zowcrIHuLRZvF
ztYLEVdlTGpavbGYk6ugQH4ukLxZatnpUB8rQDhg85tsmtTVUqCRnGdQrmptkRtFdgUMSU+bAznb
Dc2R74E6MH7ysHBgfi58wOGV2CHmWmNZVqQ4o+nHCzGLK9lwYuiV5zCSSpmx+ByxORkhmho/3y+7
bE1rDZC8mtudyuWXqRGE+Dvzg+GJf84Oc1EWADy6v26+2Hs1TD2XlCddhi7z0Go5zzVE2MDxqsFl
vkxkx9RScFdrwtZoE45Vb5zbYC3xB1CI+IwHZ5XuJwzNyy/9n6IupWANJ23DrRxf95Ar52JUUdwq
8EnX3th4ONmyGpkxvDUJXdyolP60sMTZqHWNtZiv690XBtjO9TC0M3HBxxC++OLZIJaTknbuzGbv
PQAj7ISNAEC6IY7rfMZg31YSHyJNz4MMPS3KRtS+XXl3URdM1liB/RAmT4twYCTdkrypHDIhwqJl
9atwiTGwAO3gJcPQ+2eEg+00bP3Ae0m1B2x7U7fTg1Uo+9sqr4quJkfK2rggKDXS4Jp8X6cKw2ZD
oanrQXT9Z7fXYKth3pHlQLvhgNtd9paw0eMfXhTfXrgRjEP7VGFdit5sKToN4kW91jABime58nNb
U7Uwtpqf44mE4XUbRw+fekkSLyFE7emOr0rieiCWsSPF5NFqV6Mzk/uY/An+Y2bAEihBZ4P5MvEx
B//EHMxwj959aXaAA6CSN4i3rsNRT6eJj1VDLkTQaYfbQ3p41eQEmovlCs2f86zgoZj8GI/0yfgE
S9pUpgI+xDLcy8uMPPtE3TKVG1oQkbp6yv1I9bGhTgNNwm5EENxOksTVZkHMqaFxF2tbfWmjjBfx
my1QcX8OGC05hPrTpKq+o0fOyrfwQ/TkkHIWK68OlnYdOs+HZxGFKBnL87AOz0J8zQrkVFs5zZ/u
oVTHKPrFYGYZJaswjRgZtDH+DG+Qy70cF3pzHGj1NvBYb57wMRpvmrHGEyet7HcGqWJ0/VfzinM+
li/RqV1vxt1ewCBPS3S+xPCu3hDcw1hJ5ykFSSrX+KkCrc2Wp3jGsRm4ufue4eZ5tjNdguLnQH3L
JMzlofE29gIF28jB/Im/pjif5Mk/x/KJxwi+fyO/SVNONA6FbDRcoXknQuNy9PwllkJBQdVbsOFT
p8kTp45Hlgy/bDRImlFgtP+ZO1GHvT7zqqpCkOYWBuWZql7peXMSBA0nVecRUfeTEFPaC7oTQryW
tB5Qtms4G41f99GaAXsQ/t9idvvWSrpaU6uKwZbQ1YBCH74n2hc7fOE0myqqB3VCrs9YIVRS1hPb
q1l5dOSmonjCjM/OF8/SW3yO5flFMJ4GN40YNKSFyqWlErY47Jlw7O9IoKph12mP6Ixh4iDB31TF
smWiCzqbJlM/dX5lgntUwqs1QsG0cJNMPrzNBloRhugW7s8YzAQRcxNmJ0wqVlBzUh33WR4KGTpJ
CF8fqoDTfJ6jYr0J3mpFJDusuA9tG6xUrTlVod+EiIR5j5s7EUZSNMwDHGVC/cJWXPbQdzBbvfCt
6kM69STJ56jBtyalUkWwr6RLie8UgXpF1at7BAE2xl1dsGffHkQiRWf4pz+0fIh2uAB3VhGdj4pV
Rp1zZPyygnrC4ZtHcFkYA016r12Scr7VMN6iTq2FhZf518iPKBW+nQEYI9DuOGODXUa8e0NATX51
Ortl/BdDAGQPbJXnbXHHTGlavF9stlfPid1dK0PWHeeNlrIbl95TkkMIMhX98ZVY3mUP+Vz9TfFS
9Kf5m9Emu4o+5GMw0w/FQIk5Vpf+jm2vaXFhcIM39FB+2cBNwdgmwFv5aig7rMQGA1eMZUSyD7ai
wMrHY96cMSNnFfFgd39j6TpaNayv+P/pbvJwRLibrboyBUxWl20A5SjHWrxc5yWVzXX0jF4fTfRb
OeeCP3AjcKRzRrpBsYw2idHwJ7nVHo/R00+5SMMzSnkERGIPsFRKNpdt8+yLDGwf1nyaarkhaqKi
Qs3zcJ9YNFFPzDcEyxWOZWaSgdY4XdYnQoBmXMm25N7kaw7KQCDY/AjX4WPggVGtn2h0lLrsJ5hE
k+eDkaVg7jB0hGaX6gXT05M9Knt8J0ghFHLjePpOROGkfgqClHGWIULyzo6D7aUsv9OwGL2hSbCv
GR+xzYaSCrWRbTTnsi+LFb/l2upHwnaE2VgD1RQ+CdLpk0FSu99IO7bOEmoV9KWUSj2wqWxHFgoy
UxZktgbr3aPxeIikVbsJ338NLWMH2U+hU7b8HglkYO5RXjSaR/cL9FqwSB7srFA3WVN/WsGqOdRX
9h4D12IiA5PH9H6jsktai6EBQ+j9cbfA0Wet6GMXBu8OndV01StduHPdOt0NMWOX6nZ+Sh8fgTK2
ZWZCql9iKPHQWq9t+d3cIF9MxtIFhPsCnxXD12fYIZz+EP2Xen7W6DKSYdBrybplQcTSPGWzcv6H
Qg0MR3K95saVvSm2MyJVJ36Bc3GnL7OO1RWrtRU+r/rRybs1vCUq80mKTM2Mfe7aL81OpaNCf3Zt
H6ENEw3VhpzxP0+l/9/o4bjeA3eQtSWm7Otou8Mh+cyagYFD2TgOYTYrveuSQAGHiPt2w5X94L6r
ag1SZTiu8jBHjhXXDh2Q9EVZYfoSOt/cu66RFv5LDsx9xqbZ+Vv5/Ha20rD6/pUkrOglN5Wsk5+4
nyEHzZqzKq1ATgHaJrrRNtc+GQbfvOOyb/GQ6N+kREqxWsDcnbxxPlwbqUFlEtBFvn7ONf2EkpJC
CLDSVGQQWQR9Z+jSRNvhkL5PmAarItSU+J+q9IJUTiB4o3OiMiIQ9PAOG7/NsZMUGW2VYTzkCTbB
OVar/Ijv7E6rV+NcBchCV2IauAUmRw2mKk1+dvJJcPtmrhGYzxCSFeF3GyMJzTFQlo1M+HZOTjcJ
Aqn9bSujmU2X1tnU0pLIP/KFVYhomsU5gFUBJr7GcvKRWudvRZHB/AMeyA/JUBn28JtOjsOVjjpg
MBrSCQ1dT0/kV885noYkCEyva4k72QYE84iVykJ8wruUqWJIGc2b+SW7KSOyFwn0wXIDkfN7fo/X
pfJTUQwr9E0WTTpwNITyFCQWxQBPXqKxgbcCqRJeZh6jNMezdz0wMiy9MkNjvCHXi9uLYtDNwCuO
XVfmwhXlWSPZsFmj2leqBmI+4/GxdhM3vW+9gofbFEoZlm4r5oKPF7fE33jiT1Jm3yTKkVoafcjd
Sr3XPNsX/gGWlw61iePRtg3XTzFbV6XW6p/adyW86J7ecRgIuLA65molyhQyklY/FSNs9GbjDv5E
2bXkMPJ6XJOg6HdgLwsF4lK0JC3xjImmcsGMIt3Y1wJRJ4RElUVX2WOFxdsMla7bCTW081gCHYzM
6fSvHS2Ez9LJ6X7fyVTh9xVGjZvhHnwwkVc+zaBtZs61YnKeVsolOCuVJqCp9FOKweh/c5mn6x+F
xaxhTIoJTIfIQG6L4uvzNifL3YnRDSpdX5OfF4S9Uwh6+n/P1TLupdoWM0a6wOl+9idr0yqhTL55
MIyLDFLOyJZkoo6HCvW+9FtH3vCmprkn/Ykl3v9esWMih6j0UFOM+Qh1qNXPUawb1DJl6g8ZB4Yj
tLXrziPDRHEDh9ZYm4WGMEtGzJ2jiaZTCsY61BPJl8mnTGynX5HEF1EiDkQ4WorEDV6Gvq2wMEKg
tFUPnEOgFLPio/dwoLu4qA+FgCIYkkQFQ7vtmTsFglWJmWk0cK/NUa9tZBCFHKtw3PV6oqh9PvYU
Eo1cnTzBvUFQfobMEvxf0c1uElgh+sSu9HjfgsbkZPRLJrd+GYcJlcaIxGDuDl/pM9DEFbPc07QR
BMQti54nfgf9IyalnueMCBgZmrzBKnG7f87FG1pXnrHeEE48J7m0HznQ31rB6vWRh/8IgARVS3w5
nEEFfW6AAwEJXjG0PZerkSU10EhAznuG4oKvvAEaoyVTrM0US0Wb1S8VcPiLQzIIL/BiiAFAN5bL
sr7yfWblXrdMhFgVwwaO4F6V11qdb5zBudCv6yLndVzTWlN7wKwZzhT9pz8FENaSsYbFO2KdUyYl
EX0545XQ29wPeq5dn5olU09/02pOcDYpLIdfkqhl3DB0dmlv1tkutWd6DP1eXn81CXBaRzxX0p2y
S/jUa3FIOEEMy5WU+mGjuTCYiaiewTFkQWjhPAkUJR3wobtGPEI/Y/c0SS3NeM0nzLGBDPsvy2h1
gKXhFo3UkFdlxSuaF/Il+O+XfBnsM9M4LlG/yZ4O8/3Vqduq6osYIJMRq7NtEaxSYDR/AcdnzcgN
7XA9a524lUlrkOGJTgDDyHvVctCtjXMdP4tanGgBDGN4IaJR1BYXLtsGp/4mIRi0Mp+zczgphJ/a
RB9OubBL1SaePgIh9HtH/9LBpkPIQhAjZwZpTbSajMrSVpmhFOMdi76tjsT8K4MlqXJN/LLhRezm
MiFFbZx8YljWBGVXG/WBl/oO1UQJDZFym5k4TEtGX/JE48L4TgHjJzI1utfyVKnLSo7BiEHs8iBg
HgK0ef2A59hQTr117pA2TFOdidYvJEzI75RXeTefoWNtJJeQt5t9BfP1M6xCmKO568f1ZJNXhArh
7O+3OkZhX+jRwnW7DsUBm8wKzEjWKngSrvu/fpjw/+xUCYpI0wK2JOO2ryVvbdaxuHAWD9+b3QEJ
jqtsIIHAC/X28meMo9EzMO0e4A1AuPlv9attwUppJca/ylVpJZMwhq4aFIHCSsaW/l2ccwjJzBzd
GM2iMC4ScZFz00d0O6clg+6YdzwWIPyTVfg624okU9kEDy0SbQvsInGD7OFxZt4MRLTHsuEdhOtv
yOwn7ujYN7i9we/eNVR2gvRNoBkrbEIni9NquAiIM9kSrtXOUw4fLE9T+R98JoT5bQCAO8zbCjpQ
3lI5IQx9cA3INIG4YrObXt3BGgfjWKocbXfa4loQpZhhNHSwLXoHEfNY4/Hc1Py5FvEokOV7VF0p
oqkkGJpIwZbOus8eGQTqN25W6CKm0e5YFyNEv37Bz0iXpDtNw+5OpU9g9MSijGty2cr5p6JjFYmS
pp+CGpA/pRU7x5AABQ2fBRZLriBMVwKmhgxzYjGMSjv0g20JouUq0+/PGoqq/L7Ecmu1LhnpWxcA
e3Q0vPxRBUlmp/bbL7vvFttnsgKbNlHPtwQ7Ddu8a4oFjrsGUsEZuCvP+IQeLBNiQOOV/ZLvmH/X
6RO/cNf6Irt/M2D5QanWwFWiytfZbvcTP96GurnBzT07KceJ3ZMMgfWYIxnl9gHvX8yX/CqTbHSz
amQSdnYobmhkHOuolE6vOeJRi2GYh7KfnGDA5Nh6ED5spOqqmsv+dR2yo4ALcE9dJCmCOTNaMbfu
S2GSzQLqeRHcht4DOUux70Tz1W4Fn9cyXIo8jqgu8k1D0hG+iDFb5ovGzzpAVanUtbxHdQy07xvQ
TDmbLFExmY3ntH36mZ7D/U/Z7QHUx8Ff+1xgZcAUaVbxZRiyMmcML7YmAHo/yvf0Y8PFw0nEJwNe
z2gKflE27KDvyqHzYldfJJ63mMM/YmTMB+2RNHGSei4qZJacsYyTrCzPTx17rmT9NvYLxEJZMTPI
abWbeAMrnjqIqJfiC74dNox6KW4L4mgRoSMq/UePMwF4Iem0IpHy/n77qo/NUbCNxnadBcGC2HGR
v6b28roveKCZ0pQ4xhl58dOl6Z8LoG4TIcGTsPIQYmqEe5mqB2Mj0RyFJZd05ssBe5JRcvDV08qO
q5welTI/cVAdYq4waUYeTVNXMau2sXg1cIr8Pi2g6AE0lRUf1FdcEjmE2ozwxSvZYtutO6fVKkAt
Sn7DUzpy621P5i1fT7ajpX3VgtZs+2yrKGFaAJ+3fgCQn2e0taPDFaHaZy46cGiPJLtaGjb0y1+W
o6JR77MNmFK5yoRNCdEDij4GN6JfwXcp34OjzVmBWR63hlZftoFYl/RD7K8RstWgyKN9a56IpKQo
W47BxXym9Yv33E/ctim4FeZ8RdDGG+501Q4gVummH0aNlRm9wL8slDQHZ7ng9gr1Dw/4jS/6KupW
OTcuki5NFXg2tiOuBlm8UKNkyr9XwWrhsqaxvrXYTaqHy1dloyiTYBs6pLa1Brp012oNPUD6Sg+3
yJvk2fluda2+88pDInSST/zKEPmCfoxNCJ2k+h+z6GVSG30T8I/sB7bn1YTXIlfNqcTA9gBnW/Qi
eksg6hrzy19jJq37FkCTi2YfGFen+wuJ/LmPb+4Ol+BghcDDouGLXdvz0wcR3wAxrmNuy3vvy6d5
C23GsYVL1agE2ZOomDv/3jSXe78b2oTy6EhV/BJEr+UVEAcS//5u3e2ym9DtZMq5c3CcrNjsiEj5
P3qXaQ4nM+sQZwfYeO2KduJ0jt0SjoswsbB5B9ALT2IOPMYSWU7wVBx2Q6E6O1QvsasR7tlFbDt2
I1c0hBB98cyVUEEgHHbSjI9ylVsrG4w4wsMgHHRLZ6E66o4Dca6qqkew2jJxGgdmqsMhrmchN64K
YRouwkLwQcHlUd5Nj4n77Q7EhYEG9+Wb2taY8HzJhghy8PsVTSnUNzvmrOyLIy0PRMvnK90vHJlI
8v9zJ21UGjPN5rtq8XPrHBEiCIitM/lVVsSYvNjowk70G984RwoOeTIH08WkuXzsS3rY9ud3wUk+
GsRdRMLxWIC5eR2rxQCDGgcUZJJwSRh6XGjW0pzYfaKyYX7TWL7D5zlMmTHVus7lbyuFYC0Yp79g
6aTzf46w6XWEOQum0jTjCMS4tlzDHQfEym0BbJVfLvD1QNc7/h0Hv4oS25RRarRYow59zC8/DeyP
qjkfQi+7Hr2dM69mzBFQShYvNzNqZ8XYDxnUJv76jrW38rNWEeu111GcWSQfd3Li80LZNovMUbNN
sVwIoBT0Q43zWKB1WU2QN7MiY5j72bKkbKTSRwpodQxOqJZ8YZ8ucXhJwoPTp0fm2T2EHrs5aUft
1G0OAj3yNRfLwBoZ/PVFRYrKq1yhCIwM23tifeFHjQ+lS4Dypb7nhtYrfeCq8qVWeF737ef5hUF0
JIkR2x0sECsjvioyr3mYogb2J2D/0bEyvQYuJpl9J4wfxo5WoZewrD5WzYgkUwBeDfGYrybPGkGs
KBCcLm9krpmBq5EIvJ8FC9B3brwlvLXFynPg//L2pgTCYnbOcdPpdUmQfDfCuhh2+fPSX4cxWltX
8IIvfXgk4EK9jmehAv0FHUed9vaWd+QBu1rvRscu6sMWoK/NeTLnRFUma2DwHtZID8A7+81ivsgi
pMvUBvf7GctGkiCdDRL5944nZPnU0lflEsiMH/ONR1ikXsdyW9RR9n+1qM4FRclqp64iro6iAJ0X
BANLcGGvi3XsCFT6334bVlZj2dm30twmD+pzq2rdzWK44oz4B5mvMiIqvYL0lbk1w1EsNgdyX9iT
+c2odi1jixa4BhX6oyAzLCbi/mImJO/t2zqRkQfVp0eum0haeLhcCUcK4nzADVWwEK6LwKh3nBv0
oIjSNS1w+0hkbzbZpk/JFa0/0e/sKNacn5WHo7N0nroVJdKvKovnkzQ1ViSpX3Fk1snxU21609mr
o3WDkUcuduMRG23qjOxuB3rc1sx0hLMrCyFFwGhCrTRXfmXpzjSoCs+Q37tW8EDAiwKoYBMieTlB
eNdUs8Qzoy2X2bicoRwSo2KkNvlRpqOOU7Kwj+cltrQqWMFBUadYGSPWFVJHB1OgL7ZGdfgqXvEN
t4bUNhwvu6y0srt4xvLcdrsaCaUMrRJLYajgGvb51YTFtc64BGRkRYHfBoKnKeatHuwmvA4UtujP
1buf23/uLsN8bDSGq0bxo4KUqHDpm927GYUXOfLuE1O+LVuM+Hw4nyGF2AaVp9zyd+o3HvCwSCrS
BLnIQSZla5LDYmrR8BmWXgIEERPs61eCI+rxvomHxIIOXZDCtg2Cgv9P+c2FAhIAmv45hRFGkiQE
frimBUuM42PZItcJmgzBatNbedgm+ABJqRCPqoIsMzxji66ERwoXFqNu/7J34V886uuB/mRquSuN
DaI8RsGNTqcI3VvBluEYSvwB7d+4cstpw7gN5XcY6WOt/km8p2MW3d9O9MWw4xm1IpNvsT9bjsOp
jM+5zLco2VQ/8fAHNHvFXZ63cB6ldT2RyoznZmb933FvyAeToWIQShFYVKMVa9ek2Z52YEpEplXi
sREKF8r+DEqYr5edBjAwLtzP8Y1QLLkIh1bYNJXoJoW5r1/Y3cnLlSyBQd9F2Bd4s6PeiJxpt6yz
ygj/z8gZFLIW3NQjK6rukR9pTZcURQEwHtpaxOY9DkCq1Am5+GbZ9kdoinhRTkCLkJplvNLN2a+D
cbPqVe1tK6r7A1CldplTG/ra2pVCNXzNmYz9stIncMF2pQ8ubs9Agp+NAhn8VjAN789QldFpzKHZ
Xr9snA0Z6BCREvybJw0T4KlKDGyDYiH9gV/0Dyn19UUJ565eTIyFTaK6EpHidgqWGYXOdYPydloq
T/H7t+ErleZ/AWsTHeWNhQ7WLxZbKj7+TmefDVQZRy65PLHBMd4EXmqvzeEPyWLRoX4DAV6HK2dq
bTQ4II0FE1ToCLd5/xOKBTBBVSZju8XGiT6HMEojHWT6Fq/wJVXOe+/kvg/aPJUusETXDYVnxeg1
IJ+iRDuP2ppZ2svRTrszvNtRwsPurwvzl8pan5jKnS8JdbOoD2heJ9PYxEMZ274Eqj3Rl2bFZMwu
UvrtCi9tgm3KROUqBU8UThsaH1T+CYuRasA6S5F804+GWkfx7CXFeqTTY7XtnY5cRiONcGAYbSjw
njs9dDGcQNeKXbHtKW465VP+ArVAYCCGeGabPzupWWwvZrP0hbk/pPPbmiRHma6M6ONKwpX8onlb
jrNWupORwZlGLjRTwG05Wu6Y1EvhbOvieJFz1By3Zq2ANKsnpfmdLCLc+LaLbVL+zzNxGFlBTAfR
jiAQa5leQ1U+2iA/fszgw1qlv1zWKLnZiitzlwl/rE2AfsdcdL4cYmvBKfHp67M2c+TSoNdo9XrB
ytRDb8FkHVMD1iFznJ1GICa+qzUAl3spoCFfjXMg00qGkwPzclq5v6Ihmh/u916AgA1ag70/W867
qAGlz4oFR2L1tA//r3vYkpldqEIv+KPw4u7kVrSF37GuZvIfsJ0a/8z9hdVCNLyk+iF8WuXL0Psa
BmedYIOGE8Gtn/Rk/nky2LvpGC/OzhQeKYboaJCaqwStq2Y7NBm9OA24/OtonJAcBMc6Il96lrkN
ynUnwdy5nLr0ZGJKloi3XwhbP5M/0Ts+exXicu8tltNo0GTO7AoLT3t4ORPEecaPOAGruZx/Q5cF
nOPytdKXLGOeL58nmyfiYgfZfOVCOOpDbvp+KxCdh5H1VVMS3YD33nDtMm39fx00OOgxHbHQjKGg
eq7cC1FRLOBPCEwn0Xmv3eNqYkOzckvQq3KYWAqjxsIMXL0WJ0A6dndinvbE/vDXgu5uQ8Zm0QQk
hx8bl5cEpeadheD5qyTZBB/QzA1KQRJKAtPj9WNSghCg+yAXpfj7IzENMKhTcDn40824RULAJqAK
CkAze5MWIDr5Y8cwPQgYy2gIe1xbJVezu10ndsuvRz1cmrDD+io5UjgMYBo31iAZ0Gi4dDCMHfk2
ARlyIZGws4w3ikKAZx9uvWM0UWS60IAgcv0GuEZZ+WhlJmXAQ6ZS/wRL72jQSzES5Fdxh/DJo1GP
JamyhzDK4tlR/bGkgeWx4FeNMocshUV3UJEXSQ4yNv6YqQ2errxDZFC+YbxroAKHgOmxiVGaXkbA
0ldlvn/XvNYSa/hFn3yO7cCQczBR30Yj4y6Oqy5kCy1QZ8hYYTP1S4Vme6h1RQbzIDgeTnvhNjCI
QGNlN71Q2gAOg5ETqKyQZwTVEz40HUBwQMX32X/YDDE6FxQFJtGcG+SL+PA/e8oP8VmpP4yPog3T
bpHGVqQsxP0FHvmA2W+WHg6NvH2+y3Bc437+R1yKs2A8UxA3ILh3UEdO4q65afpoQvwxhncp3zed
BhJCK+66eEuk+ZXbIePkrCUEAaOaBnv+5UD0uhg3rAxL4pw8ChOcTZXUHIJWjnn5Zy6FSsP+XYr9
rBQlmFoAq5p07iI505uGJo6lrDqiAwLWernHRJM7SL5+JXSStIQHgQAcHfbzB25o8vFjVRcYOsyz
91pnuuIH6+OWL/ZEZllSvWfTG/ztnM2f6a8wtU5mO39IBdjhR8RikUl1jMG+qbkT1zYxb0ePKNK9
zs1UpufPqK2XF8LA4c6J58svMfy5VLVCnFbODVuuWipwu88+/p3XdxhuIR+1E61DyagXE2o9n0WR
kqt1lmifAcTILPK/e3hTlqist1gTbUXHvaGmYnxvqM2uOUW0j8lYMj1Z6EBsOa21SLAdshGfNjXy
6v3yw7tpQTiD3bOvLmpB8b4GY5XqFBz5FIWtjr15AuTxI6DfO/jNSGl3r6jsP2a5CO9DU8MK9q0n
Xz/TA0vz54O/JJqbrH3fT68zg19alHx+JLEu787GrWdwLG5pLCk6qoCp5Imzh2u9kYOCK3GhjRCW
ldM9xR4QhlxQsglUAeJ+yr1i1kUh8QnPx6c7oaYdnfuXoq7J647ByksRiRvrvuBKA34q+Db7+X+J
jbAejFqp+jZ3P56LhiOgOplcA+G0z/KR6Zwr5t7c4TbOZoIqrPe66B6S6tidMZRiaH+znJoeHwWa
ooTBX9tLchZjCKkhUuPlwbpN9xmEi/L/LXloKzgZIUs5vpczDdJV+a+YU09Q2+Tg8ZKaHMfHTIyj
2EhxnEV3QalDbURWdceza1NuWBeehETodXndQ9oWeCiQ5JWjQCptYEpHL1rF1/h/6AUgtfKOaEz9
+LPrGB0uhBjQshIbvVRmRYm3W7KugBkV+fq7OlpBjVSwcmUpSAXjKnCVLtpj7QsxNXBnA1CvoxL7
m3B8UqT9g1uJkbl1tgmiPERRLYTm0be2n2F1iBo9SAmCcLU/T9X61ouUQlipxqs9Sri+WR8QNAPO
13essQuXKyu8ymrK9WgXRCXCqBFfkYAD4haThcHHjszkFTSWsY/ZGmsYQinH83Mu2Sk9fl9+uBkj
RepG1vbqfzv2NBMcf6XgZwyQezrghYc908pBLYVuECwaGUCGwVEEWKYd1ExXo8zujNyXMhtLUoQQ
Tf0VoTLQHlpSEj4TiTOw1z4b6y3Qy1R6R6fztfY5mZE19iJiTcZ3qM4Q48p4/sAtHupmfo5lB656
GGlHaBg0BbRmCKALqTWD42GWJNi98Bz2P6fGNJkaxMYus33e+1Cxc6oMJqFKzBSvWf/C/kSMiCCG
VkKW4wbDYD9+DzTY8bW942H8zwgyMBdRD00Vhx/cHUGrfh600M2//8aRMujvLEkk6IvQr4mrLia4
nmPLkg87guOznhLzAVmL3XZHvpNnvHEzrHI+W/iP8vVRc2GL5hexW+CP7hyV0DjLgsCeP0IhfVLG
XXZWBNsg7H1LO4KiL66oa8edXQvp7ZFcx2HJvfX1oyFDWSU46rfLffSJfTrb96ygUE7Rdmk3jfoe
nKpWlyIxY3LOZL28oXbJOpjhmMOCX3Zsq0sdSNMVugCBYO993ya3FtOkkXa2kK5ZGd5AzlTB4XSd
eX0HNLUJCJOAc6gltZvofOE2GUbXVDFMT/JmQWRnSMTV5KokT2AsK57iWGe+Qd9DIH0b2DJGTXvX
DLG111A/7EQtsgYBw04N3SSDJz7gaJpEB/79SYXogl5qFpPpVubWL+2vG0Q8kUwD6SZGJL7Oez9U
R9KEhKclUXqZoWnisztsPWBif6EdTaXWFFM6o1XW61Lmvi7Z55ebhCjp3y59lVpmDkmFISTTnah2
ebBXUM/ddcZ8cL+84xrUBuC7uTCQlIwx0G+Q2OUMcox7BeQ1mOfb036psD/L4VUUO98ENdfhpw9Z
GZsYoXBHbQUvqTNSddhu5nH0I62lo8Qe4nTcVil5BXPqsChFP8mF+7l5tJENRyLaPDaWCgbVz78r
eUpaxiJ1lxCPQ6qLmUqlhDbn9DklLZxGguCyuXeP+gattCHu1EiqjFzG8AROXoia6QN+JDfYOARE
5Mwaz1/ot3Dz/j1HSUBUxx6ta032JKk1snEK7EtyxpwLjBXcpSHN323DjzE8/rLDJ0sxtUyNj3GJ
NZDOZ7jhcvJaWSioD7WWASu1LIDzrsn6cnu83VjAVVIVlpOzbw/K7wayr/dpuKy6N1r0qxI/5pt5
EMqoYVC9vSbItTYw90Zkvi9ykR+nawrMCaBTA2H5CeqYuIizFDDOhF3+gEp+j9ghYDycv7CxA+C3
hYbtl0iW1dvxyCL8JZutZnlDcSfRZeHdukoSVfen78owjwUWrWLSKlIG1ZDA5UKOsrl3M54Rj0mV
oy4OvZFpUoSREML2BCLEHTR5nv0QQONljOeMQDRArGwPNIn6Usg6Rp8FEB+DRCQlJjpl04eTOPC5
aNOfFnil8csgu4NruUhdKfPo/E6pYCL4OdqQMUj+Shd3eDxymGoNdbrrmuvcCLpRD099rTJHXygO
oYVd/Ux/57wBUajuOOeOzYaU0f66KuWPzasfIDFBYDOcene1Jj7pIltkKZwpUG07/+9Pe1+AhkP9
pvXExeel4vPjJYMXYdmn1JUWNkDVgE4TClRtLazNhaNrecwqFSmfwLeFgt8V+RWPBuLPIjcy1Xuc
gbKDMMBn9RqumEM1mYez0iTF7meOn69zZu33MOFSklqk046+ChRn2mqdV5yPlc83ZCg+F5LWo7rd
nFsgYcB1+rtU1uHszysh1xBalct+c6Ce6GamEsyUaBTvI0oAZa6A1p/4vh6SM4wQCFdU0N5TBh86
lLS9CmvtUuq6eEdDl92AQdI0amrpy2tUFbiLZ/ZV6S8S6BGw5a+LRmqorD7TAwYHxgh3Wd+4vxVt
JSbVHd5md+AdOI7wIYM6cZyyiKNl6Q3YhzRKOyqdkhfba5oEYjYm9wpBGQ51s2TrKJzxcr95TdTY
a0CErGOiB6SOz7A6DPop/m/5GD2IydKh8fdJ3RZ1d+nCOtU2U87M+FjdLVauAX2CBel/p+1LVdFt
ZATrKGHpgVOURACSxeK76PisEqzwqIY8WDxhPhnRhsKzK/xRwWRufT2nOhIF8bGBD/GpY1eWpj54
Ohcb7R809X6YZFQT5si50/imlaClVQ9VdfbJzkwPwVOVr160pEdcSt81L2GyWKg9k20tZhLNiZON
5nFJC1ze1kztrGKHvgsQUViHzjmQmvQWfTJbxiaCkw23Ca5BWOFWsQZr0qn2vka9mfHwbomUNdBj
CFpyeWovfcyt5iYTSfH2gbBZpQr47DNkjXy/xsNQLC0Ii59HkAzKf6qrvaALPG3OuBZgV4uhCuUU
SSBPBCmJQie25qtZ5HFrrRPqk7FRPpvlobC5g/GkzOfDbmtruRkf/1bECmZ26tHoI8sXkpLyzGP1
uK59W4tn6uvzWAwseZD0Hl4UlTtnQygi3qfFGTInfbk721PvOSXxq1KaP8IxlITQj52+r5Vrke+W
i8QiqmbyzkLhWHbUe+Cq6X35hMsM5BBD3I5MhheaCUJJuVg9MUNEVKx0rBngh5vlAyd0sn7jTpLZ
qvregOtM87PZjjy0ezyVygeGbyvy8nL2HPm9K9rfF+cU62aWyCUckJUj2MSxUMosYEWvGWZwNh4T
wJYOoqyO4bjElAeq70iQScHdGTKAxj4AoFt3sGBwAvH8yRaYkmaEJkcivYcgJ81Tll0upJpeO62K
TGnfYPQTA0J1VS9aEXpHqKEOUk97Jidlbygh7HAqqFueE+WUEuBHR4c+gcpAM9zGpJKF45g5tq87
lE7apaPGG8OUkvqbB/Tu/2Y1feJ2dqxc4nDwAcqC45jeBqkbFiBDIJi21uoHD9JLW7+3UBKAcVpA
VJu/r3fVtniBk+vHUJZtwmryYWPntfi3S9UTs7lF/8skyXSl959Qb6mREFQjXq8PzWQofoKFowod
qIqHhB5uD1A5oKN8fgap30Vz7+cJBL+iLq1XVbvn7FyyICyaWiWU8RG1gWYr+qzeOiaN88EKgXrl
R4Iqqw946PatkWj4FZZegdevNO3LEQEfpq3vNGxcVxnLtJ1j6RCq1Sl6HV6P1P98Qc9qkxL0l0CG
sGkkHkpddebx+P1Zm2csu+zorjhjkhLnPOBv3fvfczoDsfJKmXXizwLabNW8SGYY/uldd5/iRTDS
cJcR4PS5xfmOCPuTkadd4HVzDIgjvEfFDuhahSQ4dsXAPYWtQInDp19xncClEtCObIl7ZMBmOdJc
socYjwUipCW/A7XUSRswbIA9a5+/LHtXgaX5E4FR2W1iwX4fudACRwtiYkjmlLxpTLAoXHJgLSwb
MW25Tm8J4gQFGx52cz2gBTL3GxXoQOAmqGb3rPLTnQ01LpLyuy4Icka3pC4hh7PcxRZuavY0fpMq
1dCylor9hU/wq9hIpWcHc017x9IjJDKAfZx5wLztJQSHz2JZ5FA6+MXd4DdQgzDgVNHjNUh+dHP6
EgFH/FM9z754DAJqx9iq1ebUCRHIWzQQ4cXPqpSFzeRnlnpC+vGkPcGURoaMXwwn6oEFFPk9Orn2
rLWuYKqvwxggTdxtJ8Sazsg/QqEI6DQOKFOvob5t+qiC7ttaKEIE6aYFzaGw1eHS2R7EXEsl1GC1
voZTsa4/624HOTAORfd6oIXwxxNMUAxCMGDscmps7jkSald8/TiLY4+9roV/yaBx6t78r+wbAhT1
vsYYCWwtp9t6qNVeYGZVTyrhBbo+ajgW68cLw+EQxDlNyNcR+JTHKJjxZq57ItaVVF/QeAl0BPiF
ui950nHFXb4sX2Q3JdYVdJWqJOVtzFWH7CSzCZixidmDx/p86J5Fm+mry+CU4kTwjY83A8hxfHOV
UXudhTqfbR00Jd+b3wPOHg6WEjamPSN7Q3hASasLwqJ2EJrupmSUjvpiXIhne4DRU1B0eYmL4Ty8
/dpPMJpjQ0E6eAWqY6dXVpMSaTOlLd4SCnJlFF3GuslC1GAs//3Vk9Oa6bHNn7mCquDS+F+4hpD6
+iepfggyq7o4Ap59TIS4DDxL3RlXJI2kQSTf+skZ6JLJ5eiUmUEM4cJKF+/Gz2fBDrsT5KT5AAom
eYlR2R6RS42duqk6aWvHKD2NvnDG/2NMCsIvHHg99LWDg5zt+ISbTKkOxcE7mne8zClPximh8a8O
FNg3u9pi1uLpNc3rLC/+zA3R+gdhsEfFSEP8cIIVXQEhY4HWwXqPTegiTMnOeIEE/o9WwMufT7nz
C0Tqxz1ADAK+lYYjdShXMAGykYi952WIzlbD0LuPemRIdfWCacTrFubshR4I+dElxVSIeW/l3UGL
Tv6M8D9Sq944bBlmsM65/fRmqlBcldtZ7WRxK5UvCsV+D5YA4KKFJQoIU0t2WY7cg/T3EDS2nayY
o3ff7saeB7Gw8/rjCEy9+JwVmxkbJC1f0pnJWo33mvuoKOj8k1gvMyRgkKfMWYr7zm/tUapB4bWw
BfKKIGzlrke3lFM+ur+sY2kQlyEy+TqBzIT/xdz7cYlRZ/HXlTocKBvwacqUIJ3GkOkBXpp9Jzjh
XNB1BsBdq5asXSjVG3JhhvlWCf+1+JDHMx0pIp0QKCG6oG7JdW0Jg/J4sNowHMOCNtoLO9VCq8uW
5gacqSlNchKKfXBFHoW0tKcdM9qRbpVix4TkCt2c0XX++D9/WjCCTEh50C+9IZne9E2288eKrnRQ
Q9+vWEmXIN0y314N0sIgAiSzlW2gj5/jTj42WVGRmmdgntVfqJOGo7X+3gfoITlaYF8HiFolcuoI
XKQKZlIW2HakvO9WNmWHWeAyAYLd0XxZ5ZG1Q47edLQOrJGWR+gVb23x6i+tEYziR7acgtNcObPM
7NSdLoYZaML114Bdyfb173EtGQfURP6m8BrbORBF77s+NyJI8joHLLmFlcbrn1usXQIJRAeK9MTo
Htb5qncEq4DUwmJDuoycfVFRepUupOgY8bmjwDPYjyVdZnkZU4YEsA1+Nftw0e4ldIl93KQkKd6h
XI0kjzbqDwx2osaMrTmV8ThXdTL8Au01R4vWf2m+fD/SqYyi9NyMtgSVkKXwvpe/j9/m83R3ZBLf
zOiFXEhVQQTijDo/mqVx6L9jmERm8KO8h//XcrCeATQjbJBVRkckysJAlxnhOo6xtsoYw7Gox4es
dsuxvfFkluGjP9yi09FHc1qhNznOoxmwVhOVZ9d3/1feONslWV+JaiwIrVkgN3Ae5gjesnMBcifx
Q/4aBOd5vaEsmfgt/v8PgTgmOo2ScuErKNEtvd4h3j1mJCq/a4bx2oBRHZcn9VRYtd8g6CH4jkLs
8543oJ4yKWHCnHKbCgwuoAdmWq5T7GASriZP1VKr8oAhM792GOdLeWQok/LvOt5+nA0xUrm4Py6X
v0emTgzmmgJu6w9SAzEuIASXn9DkMb2r35wnct77GgIJFxjPuLa9P5/YFz+++gtFaljXajLkoeFj
Rs4lLGo4+E8NcMowcBpZKXdIj9mX95vHD+Nc0KLC+i3LVD3mbHHXNxd/bIUGTrEAS3EB7ikNuzSA
Lh1jYQA3TwZDa9whcAQo5/blEIcD32SUVBS9LH7LScJzz0EaFAJEdml4RkYAs1InsBIClUlO2Ydq
sDls9qPkb+FknydSrSK8aOP3Gh0m8ou8xz4N6HygcjDVgweCv0ACDAeu3QHmjdqLW+9NbJFDBFpx
ceqBEJmKrXivlCGKSf5vULDB41dFQIfojii8EJJprMkLgSjNrAPYuGGusB0fH2EGl0OQ4CexJmTE
Xl31VTlU6tdFT2eomISHovRmxNmfKL9mBEGl+zvJnAsMtVCmW4zB+axbscmzR413ZxetIY/q6ZhV
J0Gj2QhPnSLDYu5aJilvPZ5lwPxmJtZ0DBWs5/iNMMPKqbqoNIwGlSc1P2eQnq4facc70VVtwIh/
f9ARTVqy5gdxIoCx6fGaq0bAFXgVtx/0EwaatzNLFl797IphMvfgO9MUqrmY9t7VUH9rowuxts2S
Cl8o3S6wI48oH9XQjyMdygY59iZaggusXcURq1Oa82v65iMaZa93NaLmyHrleGh7iCRp5y+pTCru
ajpkReuBJm/zLbCI7Ndjf0BO4sZs5cMeldBx2mrlVFLNDKO2ucgL/32NBzgLQeGS7HYqaF6SB3Gd
ALQ0XtPU0kuhzD4vD2u1iW4M+FDauhHbnC+G1IiFxq2baQVJ3SRXUfxc96jdPgT9JFlT0/YU5zBI
3WHfIpQQw0Jb5CbFB4qazhJotxBdME/4nhF91IOZHb5vlydizmN+7jweGMItraY9YtExqVvjpyv+
U/QhJQxq5rSPcFl9P0i3gnmNQLNCzPKG91T1wPFTKTtRTO1Qi5q9TvFg7q1nKFWDPfNLcUaModeR
actLgq7Xfgu7HzhOaxkkvmmKx+0j+9pu5mQtin3dMTns5q1KbcWOx+2sAeFnv+9y6tI8/6G5kPEr
TMW9G0AqJ6QcP9RICMZPz+7kpAhXEF2od0OETXUp0R8mBY7qajTYL2Thu3AxISPrRbHdD1vVjtHh
aob6RjmHMq0iR47kEF2ivPl0tAQuVkkNBNpzwzuvmb0m2SXLD9vXaBfhd6YShJIBE0cYVouQM944
9ytULiPxnUl1WrRj3do8wIZ3P4Udqt0g9+wZ1JRIFj8vxYCP3/enJ8GUof9OjQphCdvUBOu2zsTA
weW3xoLhED9maVoKf9LDMl28rRfuL0WwRrePDo337A/UhOCFQDkl2fUe+jkD3L/1qc/ybnKgEH+q
jYuLEqugjQiYubzqGPckTe9dWumINO8Hth14pQhfQq9BDVD3TI6BZgPcU7OuZmIxGXXNpODn1o0b
1H26QfdpkxbBAY2NO0nSAZ11fjLgi8I5xDjvkVPpmqjhBgE3zXN3DeJB6KZpp8ZXnjEWmb5VTz87
neQNan9GCULoiYvZJGB5xrEGQxfeXRvv4pxMlPSIIdk9j7HhMSgOAXIWCWNatkwFDAjx6h1cLKH5
M4z6s/DC0QF2qfzjBy5h4YbSMP4Hzlg4rA4eogYXhX6et0aTpOY+g8xd/Du+6ViNoActM447h8FP
vKJuar3aIRm4x+sbrVHwohqsBgsGodFS6oramqSmWky0qoxniJLF/2wEpmZagj9DztdcCPgqp99s
cEHFEud2PNjYpovWloGmYy+/nQMUtutmlSIGf52TUv97G68fOcDWC1baUI+v8kwyPru02rj33NeM
gHuDBStkHVcyIh7BIloHYxh5HA08IV9z+6thLZ/bwgVGu6GqOW0csSbv/NBiAc0DmxwN1Bj2JQd8
gGw9vK8woJXWj2GuU9/PKBMx7e4j84N0sDEcpA/MnQXp9QBOiTkwXlMpIVPrSdC5hyAuppFNJHX9
BJftPoUoBEsC/5hlFb8dBgXwKHVVRxWMO5uHyMo9H1fhnCONpU8bO3qYapzx2xMCJtqSV3L+pw9+
cPCu2ux72tLvq6HLGBnwI+jW/CiDZHnrapLPKCjgNRDv7uQAj1tfFBBUbrA2efBgz001GH9F3k9S
Ywg0Cch1+EaNxIvJq+3m3W4qZuz3ModRe5bkYEBHFlc9Pb/R2H5Obzli4LoSL+w4TWVJAfFi5zpg
jI/mvZTyGowLlbpp2XSqW12OHAa2LwjNs+I7YDKKAU/t6Qb2qLgQX7od4N8abSO/9R85YjiCPI/Q
29YFFyecXie38xV1fQGTjBfrJtNlsABs4Hu8ja9BnvIqFdKNZU9hrEZFepfLeRCpH84me0olPNJN
5KlQJLph9PNNcX1Umj24ScvkkiJ8GkX6SMqxcI7NSpT5vmZ50fWTAwBbrvILIioNooumjtD2ZhHb
ew/kIHTWZ4TmuJGJ4P8s06eAS5U7tI3aghS6EbZqcw469/Qio9QmPRoYS5oor3yQ+dQlcXE4Momq
H4qM13ymYGQqDrW6Q7PIlaZdZ4r3DfAKC5KIb1GKPEofM8Gdfc+4eFj+9dWfHeE8eWCG6nbq8lrR
9EOGTLuClP0pnmKmEGxOXtU6kf1+1e9eHhBtKk9rV+Qdrv1EM7BD+5rHj5w8EYdJRLfkQ6m2lzP9
gq+E0Mi5b35inGR50I3QNJOR0/uATtu7lxu1z270CH/0KWaq+R1aXZ2EOhNkakSK2cvX79Xooc5t
Ei2nTU5uAgZeHNIBbQyWbPLHrBcs+XILbkF3Y4ct7mbV5TCCfG90RZInzt9emzghyQw2gO3wk0He
BZ3osSuitRli7AML72Oa0it2n4XX4PAxtQZHnxWOUJVMiCw4FgyhTrrPn7k6tm0DtJuL6g2UQ43/
7yTcQtgYv9NDW+XlaxWh/pfIFxMSAE3VsruEGGkwU+UlHS/ZZAWRMIvnCrurFGGAKmTXCn61HRxS
HuhhZl/z/QdMoLw/tenx/VCMH3zlCKcduPlTmONU1crYzX5c8G4w7QaUTbdbMOMtMqTSvNCeeXMN
GbAuXN1jNTHHg4NU6K21/lqtMOGHRHcG1PbToMiAcHUWtREYmgRKQ2fE3Uxp+1VBGflX+OjSc05F
BgM2JTWl5l5KLyeoc23s/3PRX+JJgSh0rFKWCj3RntT2bkpO3tCu99c/LjeEGlAMcl1J67v1/Iyv
wTMGYH7idCpdSJwjZWYHE436XfAqslZxaAG1yl1QjUOwyQydT2lvV6G56ZoO0cw0W/Wu0Of9S6U8
RcEYwZaF0RocwB9Du1lWWS32Kozyvjtn9a2BuQQA165ybWogEMSyjqkz3yl7Lkui/D5fq7O5WzF8
gnjFWOITXeiImo2nIub2r/Zn46dYftqeFJqxi5uI5oEAmqnhyxi2+W4FaALIxh3btKhTCh0WEpi4
WKnqV/DwGJon6j98q5F6TVLZubD8goj1jgezXckOVgMY7rg2EK/VVvkHhjr+p6eKtdkqV2Ti+ykB
Xj2D+I1IrzMRbjqbKiowL4c3TRHwnP3UZ9ow4unZHJLvmzUeoX2edoy2V7CtQKE9qbrYrsmUPepr
gYdwkQkeAFgicRg4g/vaDWNJkRsJ1ZZc7VrjK3u1NDdLjzpRhXlPXbY9ypXRXamHgcwIKQ0ceEtq
pfTCMagM1PZrZozsPhQVIcwE/XXtYRslFAII68WpDeegIKpMb7mxzuPnQ7LptPD6aP9lydTXQfV4
qWl8iOlfgyE7emOF/fjAEqK1Ktm/tzb5G7oso0Aa37j0CsvUyl7rUVqnCKMIFCPlMXQQ2QgwPqJy
jTfbdbu3ywuipBEhQDw8GaLSAfYwJjF/7biWXUqvTGWF3CY4jFq+449PRFhsjAuFMkgR5vphqLEm
9YjnoCBEcBgZgMMec5czil+ZipecHJbqDR6KkRSzyg8Sjbn5sZ/z5Kr8qORRoRsipiV3YBDaEcCH
U8jatiBBRBMSvKMAYiOr2CdnzUDHBAwpG2D0stely3/UJ7xhsYtEFnMD83818n0dxK8Qwk5LJ1g1
YAW0MHOhcXh4dybmewYXel/CVNUrfXATC8SYFg864yAQEfipKz/FqybgfbIGxaXiUZtmPoK0Hi6b
ZrzR0wqIAl3zPgJ1BLFHW2LyR3Wydx9aCXe5TivQhSQsEjlwZJhKszdn2mxMvJJ98LsgEC5JNc5s
FgV/Uq4T4hhwkWPn+laMljDEua0SobC/xG2aiF1luadlrntxVqZFdpn2R65YTRAbe2G+C4jZLd/J
CqHG9OrQGp3G3S8pPBip4/YsUA8X8qu5q8fAF/ICw7L+UKlCM1hcIkqfe2wEnD3K0w0RSHKrDYOb
2K5GGrsg7Us6JWslbGMpJHIitOPL8nbeRri7VatUYJ/nPfLYlbwW9WxNuP0x40JNodezdWC7hABC
SGZJ6IPC8GlgYnp+FbdOMJFC2E8mKVEDwS72jRvqahWgAigVaSjNNy7IsDcqzbee8nUHvylpjVM3
ErBxZyyIUcTblaHCxfB9RClNDLhfG/fbwDkMc4dT/ihQsqdnXn3wz6UJxozyrDPWiX+n0LfCRPUZ
0NsTmhWVOFp+VtdJxT7mUP/btzqDCXMhRkbHTC8wkPxJwbxMnJDG8zzQoKMaa3Ou/wmcJaoDSUVd
gyBk9FmYTCzDtWsmTenqA0AwxlWxVfIuXhvuN9X/n8RlLcYNDvzAVvwaiylySNlyimf+QyZJaMZj
2cazFrhBT9eUi1873Nb9NO/HLnMtn3YkoY9AXRTjcjlVu5wXvOd8QsEPDUbJUqjEdjZsv4xhoPPk
F3d84/3loa9EpVE93fxdcAVPYVWcqoQ2UGWkfpL3Tr/PgmWgpahs41/2wScOXeTf46geDYuAnSTN
soRJXYs7DdWTSzZWvQwJpHBYM3Rp1LwG0ysjdE79rUs2zGudy3ff02fODVFcMffVA2RoMK0pfAvg
6W7hpxFnk64kaqztguxKN1k5XzBSfL1GTtjycbLswguYQarA/S5OOKriZOXvXPb3myOWWEGaboR3
eHsKpgptkvvONlbcPaYuLz1wJtrL2KD8y3Qf+HPzgrQxrDtiRrANIsdyQuEInBH+szcMk3rRRVwn
HiAtepQ0XTpasfYBQQwlpP7J60lP8S1O1XlHyFMHqnVTNz+9B87Zx3AZpZbzefxMzXbdb9lcJW+x
J3sy5LNo3EReUWvPF3UY7t1dmO3ctMEAcaamz82nbAkyJHA/Dtkemi/n+2Yq8/rY0W+eHDb2+dy+
sbEolaWBLKJ4Tx9XVDpDL5BrbYh08+nFtz8MIwujD8Lx/otCla7PLZ9BbQYHiQ5VcQIqfjwpz/kZ
i7L/O/TK8LxzhbbfCwM0CUItFC0MyZhPlzAFWyjOBNlfr++rwUtXMwwiKILvG8JtzoLXw5Wv1laE
fZregXVyg//5HEdulIueumSmyKQE14BlLl82VZKvfG2uiETd4bDfdZZ7uk4IXdRiQZm9mQu41KQp
Cg/WFnJj+pN5TParJcWYgQCiwD/CXhuivSbhCtuDhVVKSXH3ksyT3EPY9kKqH4Dh3F1xb9uySSmu
F9LkY2h06TwpS4/hfyURu3+TNBoWZqsIX+fY0XMVwUeWrOioU5brIKmUhTJ+WpuVTqG59nJCoLqp
tXeHLwLzsrud1DJr7JMwPkA2XEtskDApWbn6QZ6zXvCmToj6NN7ocR7bF70Myy5D1y9RQdCVETiP
JkipP8p+KCJ0TDxsCp52++z8PkKWP/ZCaK/VIO7mi0/3ZsfAgFQh1FhQ4QYYPAGM5/xNfgZg77uA
Ni1yTIDjqlL045F8sGo5SofrDftyXb/WiT1B3IeH/HM36Ms99h5HRl9Y18M0zBOTWx4X+HFjzhKQ
LmPndIfcmSmghwOQN8f43mUHOhiC+utZ9Y34gJ5IaTBwInXgo2SAzhsd6xRDNW7SyUG6dDuuQ5C0
Yp9ibQQAmTj6DS/+CpUp8+lgKlqXgox5eV3Bi9y2Q9WYs8b+WZ7f1fg3foLJCdwZpvjStfCtBb0d
7qNfBckxfH6P50fYuREfHBXMiutguMmN+02KVzw4Zt3OWMDFIlF9NknaEZbJxgsO+sC35X/32/Fp
YUCXZRs6nBTKSKLQfazJmYn1olL5vZkssx2pXN4duZE0ug6mgr0qQM/f/YobbyXu2kc2JU3Urx8e
d0glDuvT5g8ds+dtQhOzHcmhTgf1PhEycfGTQJugO8Muf7/V5sOLZQzZt9OWhH72lvGQ+IkAt9F7
Ajp0QB9QFTd0lui/OoUSEZKVUfFP4vaiXunr3V+9gEkUp071MfSDnXk5MbiLI/f2v1foV0axdryR
oICDlxAW7Ksor/WYd48f3yiWLQl87h6R1tvgP8OGQ5eKgADftNrmQk7oTR02uWZ++DQE8jh8teEU
TRj5IR8D8gc8biH9jQxP7OmugDQV2L7BgJGtdNZVD6Owdiq+Xfo9E9IbGmYjJMtTt6uNNOBb5+aH
fWOOSdzJnK13+Mpbu8TlK4OseCYvL7hcudbeCom7K2RjSOdTW5v3anZCedaXzhSQJd5EMYXIP9cL
lUV0u8iawouVoevQ2jT9WQ25gKqIXA7qFqWFspD8KvFHvK5qr/jUWtGuPxeGBDy1ocCdhnz04sVA
mJXc8JZu6hZ1PzvSUkVjJg0TC5qbp49FXL2RQgF0Ij7ZHDBjpB78ecd4jX1CxRZcpPJUXQEeSVKm
KyCoETnvUxBz8oMHR+Bsi26Qsd4ZGH5DPGj44uqE71tNz+u0o1QJNyDMgo4rCO9d/XT26zSqum69
ZGF5lepWumt1GOYt71Q+fte+O/xAHxMgFmanEIrsiEHkCu2SDQ8o5sc/waqbkL9/cPFt3uHYdt3C
EBxnv0yYUyzUS4FWynajjVjNNs6RR2ALzZRi8e6c4zjp+bYsZ1SYsshHX2mMdRUgE9NstjFjY544
/+QdiiLb0h5ApPbv6Qun8OxsgnIFPhr4AXRCw3FzDehuWabCmMaT3xgtPwDP8NsWJXgrZE0MB5vR
+YwvMS0NsnRIHdAIspVX+Vn/7a6abg7EvuvdAwnnRh1g3yG5lxiQBOXWSyy68PtbgOK6TZ3l1M0d
MCPAAJrJvHPHwVQ5o2hesqhuKZZCbcyNhFJjyLqRM7jRplMklkmj+U7Sz1xkVhJuSLt25p/k+xc5
UN9ra0zXuyHbN4P0NH1MiBu6eo/C81W2Pcc6kjFh54dSMVMmbCW/KBrFhNy7KLFSO3cIAVczZxKo
rFt+uy1ixDGkaQuj6kZBo+dUaZ4MLSkjlzIPF6Y4OnzWv+B+IFuybTPlq9lwtMy3Fuoga3i9Iaa2
X+KZ1KCN9uTVmae18RVMoIFII7bu3I6oqAQee6aXx9yoiiYU6ubnOIn2F+0Cq8fiT0UZUSVLoo1W
4PQAivpLqTx0mWzVzEcu8mMToOBDdc0CwupwoH8wY9duwsK3PlXgAo+3qhKgIPQ/+ZYPuTBW36d/
zpWb9yo0Ehb2CqJee8iVXsmRbL/jBG3WfaEz8QDEE8L4AdNDN06hEvYfaaFmmL6sSXPgY8oz3E5h
htaJwORzl022/Jj+HHlJrjuNAKQmrK4rC/a82IkH0pnRVobSCj90oaUeYiIDjpLihTxXAit3CTu+
/xsMQyp8xYoJGzeUwsmFv5GHs3eoWqvZ/outwyb5JPAX6CeTD4e0BXaeeFn6Be9XMV2jOlrUUiDC
mjMLr7h7Zrf353JbTN6KIyA0CDUTrqf/tlDyBhDk5gSJrtUTxWJx7tVIv/NVjBygX6POQWYTqlzw
r9fanMw62+SPdfS4nk3vpSDXKyPJ1UuB6uZHVhjRl1yR39Lo/0cz2AY7X9awoXNOz7dKpgsETTk9
bGZaTR2O9PWVTDyPD1q5veIy3E+bbZSdhvMyZFZrUb1SdAIQejWxa0cHgtEHcmBibEVMwAhHnmrU
jIu3OJLWHMDyMdlDRtAp+rbOezHhqPaZwZ8sOXmWRiDfT+ykbO0ey+ca8CRz6LRuTAuqcfUzEHyM
9pV/864/oYs00Ru9Ju6HbnIQaggezkMAzwMbYdHWEQU5Cq5OTtGeB2Wj2snVOloA2yKRyGr7PVCk
L8LB0p51cuXMvk22HHVzqj9KvWcarMHcvmf5HCE6wXOqKVVuLPBo840errQxBW9BNz39CIqYsPfC
GzvGxuHm+74RoFbA3/28MGNDvmEUmMoWn9FlEmMKVhpCyabpztsRHBKCodi29LpfeqvbKnphJFj7
EV78w1ZeRn1rkzQsYx3n5D+t+ov5G/MGv+DVlrvOCJSU49Gzl/wZa08UmJ8WeBRGg8UFpwDQjrK1
9QiJaN/ENLEbyB9zv8KXmwvEZgzKwM+79VAFlclDfQCF3Lm15V3mgC9bDQddGorYKI6ResSgDWts
cIAJzp16YaZEfFyX5RQ/Urw+d2jHYoWX34p7Nuw9MAj0NDPNe0smGQNebuRI2ZSfpUoU34Axo5QU
waGKhB+TPIH0GzQANLHkoAbGp5beGKyq1mYAmQluUTgYh+ylGJmSFCCTR0TvexnFYdgpFvT4nw68
K83vfTv9VLzNwb1JbPoDEcXLY4p4wX84+XZhabompDJ4bhbEuAbh+/kJ7LJUZ9XLyry6/clpict/
HtiQHrBa0GbEhM4s2JTXPWRAnp0KzFvjLtoG89Yg2kH3P7B5NdB3d5K5aq9QBHXm15GPCcxoCft5
YhMrXBXB0WZwUhLm2lq+B9tym/+q54bp3Itwc7u8MefjUsDQYD6Cbikf0VBPKK8LcTtGhy8sTdbs
Xpi80GFgNf1PHXZIyP8gLTIwAwG375oNAX2ebHATqX3midQE4nTzuaqDdG/dxYbN7UQr4gvHAPFq
siaU7/4HINU07GaxXT2IOjtBBixBTHeKVLdUtZfstyZ86looQuEEsiE7R+F/t3NSWO4p0NpHN4Lz
po2fcJk6rixPC4tUA88Nt2VSDXNBhNA8On6Xc1EFxlaDzkqO5rZAaTT7odEdKWvJhawpbFXC7xwt
hig9eikR+PI1Qi6oZXzjnqny/uUs+Kw+WYmCZCnXjVceD3GgdH6pjshV1dSHr+F9C69pPOk/kPZo
GAknkYYJwsrTajdD9ikDf9Ay+FDiD52eq8cV83EHl1MQsVGKQTL5WcVCDxEPAFrYFUrsP0mCTO3l
QHie7B/UGPJ+2RVPJXHj5AqLRsbyTozC5rjeWZn9jSAtgdBBNxbS7hymM016pus4W7m4g4oIz1yR
Bp4Co7NJEtYr2wm6exerurGAqZahV8wvtnxz/0kIWHiiyue9p3ZqF8tXG/PDNstgwGJAARRkhape
1kC25XI3jcvbFfy5El27/3tL21L6MocToB6XFjYDttdmx8mxKNGgW3oO1C44JSBu09zmP1rd1Tfa
RMvDA13MWWKf3XCFcTGVvSigM/sWQXNIDsNJyHlTdo1nVGUJgzObeOFE5OTg9gnwibWTtf5qUTk2
MPlNhapaOkldcqoid4mPoMmWQeeYt1I6rgzvbB1jui0TUA0jjumJ5x1heZQI4CFx55B8RqPRAAJi
sn61q70NwNe8V/09A9TO2PiB11yDb+0n9sWnl3RnNO5eoZ6s/jvUhF0dX+BW84GqV8DaLieQs0ls
zW/JsS/oyUd2udr7NJsj2JAMLoTf72iBO5aJP5b0QOU3UNq7BzASbTsovQbgXU8ksQpHoB609Fxx
js91QVfo/jGIwdBHOf+3JZk8+JE24r+Y0RDtGHgFJO4KoLEkIp2MHr7j+WRoxT9OwwvuCIytDI5n
FxrHv5eNRJUKOf2cTDZeGzNUZgjMzhI76iI0b3stc2FR4l9SudqPgVPiv0iAB3tAz3PMxwekYqQw
xpDC+hgXZu8VJH6cNlLma7VDQSxxbYNcLod/1YVAuRzEQnkfC3hC0VxtbpgIQPDiCEaUiBSK71sZ
LEs3mNs+1R2L8gzDHcmkXNQoGu3odb1xEQlCKgxzQxh50TkWkF2wHm9fkxwfSv1jn/aGZIrIJcFz
mKzQaJGRTIPmL8oy6wzlbwrpsinX16Lwka8Iy0ZgOt9Rwwg2cJv1QOJXt26ay1LdDsnaNMxIg/Gl
419Tie8ZcMUpmYXHsC3oVJsGaCoE/rxxUJRBGaiKSP50KXoHycepqDlE7Me2AEEQz+iivfQzWyW/
67wRi2uq9LDhmYEDZqzFaa8YSDonBc37E6CGeVKENRHclxn64IMA1KeopWx3ZW/mxnq3XbFWNsFW
xC6NLkWKBKY02IxpJG/T+gbblTqhIt2drI/elmazSXOrBqhSdCQxdrcHWHWIqXQ67OEHVIo3nznM
peI7PuIz07sLncl05YVOWR5QqiUVl5fU9uJDMu91D5/xm2wZbOQtYyAmGyAiuYRrlTGIYyKSOrJw
vY9hEZ7R0FuKFJXA4lrykvc+lmGPQnVzeLDtb/8AK/XPJDScr9umD4gRYpBNoFnfBG+Oi897yDe9
szLrPNpnAaxuiS0M/us5tn/ZAy4QhIYlfbgF/sr/HGgzdBbNOf+zNZBO662f1lWj3/xMcsT0Aty1
RkSELbXm5XOK5Kz8sfdZOgWVBfmbY9NndUy5PyoOcwGBQd4B+rocdjnoXtujPp6WC6iNvb9PkhIr
8mpaNm4lslYVcyOHNsixamU8rRDbE3M/VsBWwH08lo/fHoH/a3c3Iipw2E1P8sxmqXDFRYPCLtka
qfav7NA493M/nNijrDBX8hUVfTzk0N/TrHnTlgjJ81OuQIeXi9EGYJkYZA93ExcJkLiK9u/G8tdh
XbuXIgFWGfvMuIRW3jMcwF2uLeCsRu+PYXJyA8Tf2vz+W1cr+9SBBzyZeNbeB5pH91xZ09Tr+nW5
hJSJPeaU3V/D6AQMlOwniVZRZjb2cLpPJMheLdAnAOHttUujHwdDe8OcgoFjrIpzVcWUJJGIzYEH
K3vDbmhvHERS+jkQHtSoZ6WVD15mGBk21SSwkaOQPbrAFltz/CGOINFFRZYHyeOy/Qc86/PkLEWw
ypG2MJ2cRNpp1GVfPnwJPLqGRlbyJqhog6gMqwEW895D0JdsqIRgNMgTQvlJxfTBeInunlaj0jeW
NM0mcjCrf0vP1lHLDkfXHN7HaNQ4Ocd/WI905prfNXyxNeJz7YXyw4mDV3lXJSuv652vHLUOLxjF
F07POlIiOZvx/uS1pZnKPoOz7OFLvl3HXNVM/+tqdnNNm2Oosa/gJrDDgyAVmgeqXa0ofQe8z0Us
wIZHoBq0rM4gVHOqXtU06bRj/huS25yvwiLh31/S6/LuzK6FQdZhpHECgPvK33kigsDRvGhKPXOH
IlxxfRbc+eAiW7t7PifsOfSZ46wISEVxBpKL1oewD62C4g+NjdgxdnYrgRTk1jBJ0ubU7wBHeFSH
72z7rkF8/3JJ25PjWMZTk0b5+qR+gHG3R0DyDidqjVxQHILeB9IZ6E8CKEJpFWRwdQ4+Xe6/fP/S
3TQn88KMFJz7nE+k6SJZw2/+BeUxO0cEDut4vMZ+/skQKPA6Y710inU7JMHoZKFNBSoEI87suhCH
eM+MnlpCj0m1RDGpwRfej7Ug/aNguoSYOnpB3qlbAwcglHRI+FM53VyoUJU2XQ6TleQ2/7nbbeTy
SFl6V82NJlPSLczekHEEYclCCRcos2u/DUrQlURFVvgykIRVSiLMAf6YCeQRccZoUwQ5eMjO3pDe
9k+4l1qYN8NKg5B3y49kivS/h6dc6fmRMbkLMCC44dR5m1Hd/EWvJ0oOeW5APk64mWQ0Z1lhNjr4
C0+L+CQfqp6cwT25/dfqG0AOBvjTsO3KWJiyGKyO6DH39+xCu43ZCIw2xj5BdkzCuP0LVRFo2ks4
IkCDsJem1xeGvF+Z146eyZWiAhqiPgg9s4rJ/3ymd7cqduI9C+sA30M3CZCVFx3gXT1eZ+1wyaLI
yAY7DdOaiDxfTjCBE2LfIZzO+wSxSRL0uhj7WweyOE4wwUGrvaR6Mq8BKx85s0BmzWcL0XlX5rZt
cp8AuBJqoW1Cficcoz96kG4I9z6UrSaRxr9QZ42fOdMimohliAYRnjsc5v6NH6n/FTod/0W8+Bq2
6Rw41KR40AuQjFM8nxQlz4BZZy0504E/7cMlhSQtd8R/TonEmyQ5WejWi7Mere8xe/2Fx5a8HK1m
izgJzMVMdnZSo59llGkO9eLp6Y+HyCAhFXEA9ZIBrwXlg4PN+GrYgQm61OxXIYTC04HMH/S755Zf
NCm4Ai7yVtgZZHvkEWlpNbJMe7DHNhFm/fQtIY4rqIgzaNVzmcTHDLU7bLD4lnbBCfRcVFQDufYE
sO2yG8qQNSvQvwCUMC/9NjWm/lh6E+V1e3hTKTBLRUQhCm36ACzoBJPhepM+qM91b5sM7hdzQ/4Q
3BLUKRQ+wYydl3hl8+JMEswYW1lOOdXVpey7VJ/sKCMvoTe0VrwC2RTPBDO/WjVGi1NvqhW2UnuJ
gTWDc6LLyq6cY93ovPsQD8h97eJ+WjTdOaUC82T3cjMSsp+SDQ3DMXcKuvHQ5wNz5fl1lIrRGAru
OJ1CUXK0AxU4rK6QtSdcmmkluGVUWn1c5IE6t+fUGeRtTnxxS4eZ9iuqGLGSMWrKpKMnWC//QlVS
7jE5C/DIOLlwyXNFWnwRsaSACR8sR4hXU2VtawhhXowaLkAGpnv9TtjKkbBQNXWC2C6ZRWUGd/Nu
V3neaP2jcH40uB0xN7lddPB54SOGSXRkvwhgEJYkNuXXo7z/HG6SMXlpoRGbz2EDF+u0DNHSvN9B
6dOuTxf+7ge4hOgaYuQjILypxBi9+fMYhIM26+p+LNT5Zm4wSJVRRCfws4XobX0wS5uK2SH2bOeT
r3WiI5hEpAeUW6CVTQR/+02wCkanJOuf8fJEsns8dmYlDFctCTwt6BIxw+RSz5enqeoGTIlA20vO
k2Bw99RtrDtfu1uythMOLOyhbcJJWW4xB1n3X6bIS/PSlFXwkpTUkD+jL+2klZXQ6gwqaYUeeQkp
bgcoNcDVmDkONXuZqG1w/P1EcZL0+pHcTKcfwYl2BTlRAuCQzg6El01DZBF+Qbs15cZlfZGvYpUS
p7YmVcTGql2xE7L9nXL3IIbONNmUh+gADRx7MKBabA/w2t0Af7aUPrZ3oCZkCAGB+cZXZ7sMz4AN
Q8hjAY7E6hj74a54ULiL/SEp9XVcoUYLgdbYzyKfBlcZeEguJ4XxQkmloGPZ/ELO+zMcYWKoTDU5
Bda4dVqarr29ppVTGZR1WYjTqVIcV4k8sLTsyBa2erecWhbYE2ze7TvI8KIAp/ysRVS8Gpu7oSUs
zPSHYwYOaYXO9cPlOS8YAEfRhMdhwvqJyYca+tAMHStzEn3vQLFIKpxi33W+2am+07kNZqkNo949
fmaPvivjAvNPsY4bkSOy9F5JyooLXsOWXnRTk884u7HPFCzabr+53BWNNvY/nHjNygG+fPnBB/9Z
3J9jOP583rg3b+PvhI9HdEpHDeXp26Ln3OAnq0VjxbJVXxWDdvKPTyEBP27n0+YpE8waXWdKoPw5
f2GYWVO3JFjbTfFnhY47+lYpVFculsbJv2TZsvNxRI5CjBYBLIX72UB2o3NxgVqG9lvI6N+sObmp
wCQP+FKnIARlWe9zNbrbbEsJjN5lew2hRGhPXGMfJZ0Zm4d6BJI9sBSVIJXEOdsEtSa0KfK0Yd8q
bpv+6uPPZ337Yvn6ukLOTSgC2h5hHjPz9zwkStGaXbV6LuapFgeuuuBjWo+bu7wT1Y4QJfEysEOX
G99ckiF0A2uvzh6dofWKsvYzzfER2P630lDFNp0wANdn1eqvljoTY4WhoEXFPWAG3gr74AapznxI
WSCg0DIAGdEYw50rJDUzQRkScXcRAG+kNQJjV936zMDQ6K0+iVAvgRl/SuXQrNeo//M62d3aOcXb
hHa67CvwiUU546D2+d8GCGIcVNhpciFVm0ecxcx6vPvCMQMgStjd14Zvo8zvTgJSWvM6yyTkmdRx
GKynBbxQhJ7VfMx3lhoooyynvlP6jdVhxaeXP/8wjKXp4yrHRGZNxjbuASndjOvSAv8uUcQSdBO9
HEZ8SY+WUlxm2KDKpcW+oaPOF5v8lMriYjWqBFHeA/F/ngmhCFbesG1Fc966HiE1Eh4tOu+ql0yb
WFwHkhbPId0bT2a38pYbWdjj57XCzCZ/VwxqrdrxzUAchUTmYSrvSvIqAG98itD+/NX3RQtXQKMr
EJ5p5oJnRru9Pgvl/xucHyIgi2Z9CUZih8zmB8rIfsoryDKrYWHNdCI1G9yEn+sj5SeMZRuDFdwX
v2xUxzJ7CJTAM6Nk9inRsFkNUZxE5TkPlPKQqt4PNf4SK1tGg4rAnS9SFYNzirDoXdUVeU6mNX1Y
m6gVF7AjcP/VYSipHP35GOjsmPU5NMZqeBx7S/cSXKAH0t7M0nZc9RHcIGwH/g8PPw3gmU8AuyDE
kooFYmUVltv7J0D5GgXSBR0akkulyK+FzY7K6ELqRUv2dTgLvXlnWhN5OkWMct+X9kAvw5Q9ULBO
JUPLWP9BThCVdF6k3Fca3ZiCpHWExvUOTLHwJzVaeDU6W6JNhFIHN8k6zLfhlAvAuUGoxq4ToXdB
+wMuuIETT2EPR5dVKV6h0jGuveAGQVbCTSV8HTlQVhQJyYAk3p8hYZTo2mbwDnfHEt3fbFK75xOC
W8VGj4FHlr+aamW0lJH60lRJkmFXNkvzJ15hmXWyJD9dTdX0IJB2OlDBT02UyWVLmRCACIMNy7IE
4Lapt0AnlZ3FP9C3T3qsJ3uLbDHzlAtSMMZ0B4V/9kjEnBlBMShxcSqPiqIdc34mWiCBihe8EBpN
6twgHrPnlFWi7IHs21khg73FmL6LISFBbDxfEkisqqyTZLm30DgfBikYY+nLkAFQ3DlH25hA27Wv
QmDrG7S0fefMeRAm/MBjmBv+o2kqmA72yaceY+IwRH27IpaF1hDKSZLpuN+Twz50Z7Az2WYPAJNG
AV1RcN+TfEjE1Q+DONHsaEF2HcAMiwVk7xZZo8f0NeHOHSSwDbJQgX9VuFcxPF9nOeeNlXdxn/WC
DsydcdgPsexSAf/gSGTyGyG/XpzL20Z8x8WaLyO+Ct4vwDLOUaq0FRvOs98TlqMazBS3XzWVt8es
eKQZ/AF7tCL91mAgk3WEtZGRmuJHZt2D3BFvZSpz4CalsI22YTcgVgchx98WUeL8gduPHrhJcP2Y
wSplQSxJBU/3FY8GI1YDbIz9dnEXlWL2v31jlT6qRsoBenjOpjr4MfbyLOIHZvY75jtN8YyAIzct
D53fK2otnIEU78PnsYoptelt+E3LU1DoJEezw7WxUNQsG880L3R5VveQbqcBgoADRLOVHNEVMtPQ
euWPUi+uKK0R2ZXsBtjqUhfq50KjKHJSLXP7b9iECXDAoD1fw0870fIfRJAoyNPuG0ZvB/OGca/6
dM8dRbRrblq4O/suv3iu00iA2Meolb9f+QJq1RL5OuMe6S9uE+dOvA6eAWHzoL7pOmzJpoGp51Bn
1g67sIIwhwX3FfkTk2udylTfsraFT0jyB+W0wwjfi03gD7YqJcHFpHrDxYiDUO8F+ymw2rD9TreF
4gX/eWRG4P16N3v64a1HcTH/+sBgL04QxqIwo0o2T10hLi7ZrRr0miy+nF8C10itPRamT7oHaNYB
k1aEY4G6aZAzydJjni7mspnylmLZPPiGRo7w2D9hWRfD+uFYB8aMXKQYJ5tCCLBpU0DmifVd8Hww
gagEJPGEFSR4VayZsvDgSKCOmi0+3AUX9pdk/+O+KNGRC1MGRymAwTx/+3sDpSwZd/FEy1P1z21r
KBC3MNVMQwmV9hDlhM3EACtuauV2X7pYQiVyemTsNoMhEYj0uWbxczzBfjnTtq7jm+KrFnkmdIzk
Kc6GfNGDdx6t2YeZNLewKu/1fApPOUVYM5oknN9u1N96laEjRIPw93LuqTqg/z7WlzTHxxVJArU8
fpgMiYILWX5MThGb6EUxQED5ydRlNc6YqUUfJERMqNiUAxAbIij7i/rtLCNyj3Lxu9d7QYAHBsci
YooX+1BlcU6D/wqgHMbRHP9ykWj8JxyXvuPBbHPyMYx/yu8ZhukmAu8keDATU24U5dZnRwbwmVNM
Z/Dj21ZhH5kWgWzqP50DurJLHiORDM9GpO4xZolw8PibMKWdz3qYjSDrOfwMbPnZszqWKe6GytQG
dkwMLB6FnV7Au6IWS8klh8tFxYe/8Z+wWJ9m7e1M3lspX5o93AzpEa1B03U8kVy8rcgztiqmgrYZ
VTpNSr/ljCokbv/ciPxfVbAUqDJQ+NOoAGh6IoXojRmsyfHs7LePVtx+Yo0ZcmR/f45xlhlraJ8L
s/tL9Kp3HAksaKun1GfnlW7489vYtTbqkL5GWRVvaeOUaJCT/tARFcy2PujVDidJkTDAcnt2xjh8
o2+s78jUczHB+NGpNMTtpOgEoww5wqHY6L8sFMn1ppe2nFSn+SckHZ3eEORyJHjsSNx9GHmyC2Au
KoVWWjAgv6HQHClfQOX/V5qCBPi6oKWeAnITcF6n/SdLX58TMNs8EgTrlD19l1YWaMu8gqSrdYj9
F062z21N2Pe2xiO2FlAO7CPLLPpRecjWTvm7FqJW3E6Z0S2Mmz1EDRZXXiuO2DcpFm4i32amczO3
GW0PPFgsMfcSgd0VQcgr/0TFKSDdF4u4qgrPNOKOwnfZA0Uq1NWcmV+2M/sb4HMym4uBRDVd42P7
YOOXVWeCCXmICCa0vk4dQtndDRMf/6K0Cs0AavTQNgKps5tttVphDCsbMxx0b3m8r1hv1ui/olj9
51I8Ndct9MzTkuncPiQshjQSaukGq+8DXw7pyTiZqc1KwS6tM9MkYrNGnbsFcIU22SP9KM4WYc5+
Zo7PGLST0xyS/bE9mzgXgKT232bRXuNtaqSk8wweKMsXxdUwtLfx86RL0F3/4p6/2/YbdzQEsbjj
UywSw3ZYsysYT8aHdwlLyTt7Kx6uWgTf4r58h+LwIUwzTfgel32zRd0iUUnOTrX5szzqsEZ3FDtm
eY7mdK8gkE0MyhR6jJkjZqmllYqjuVQkCpUTaHrt6jciGVu6M0ivm3tcs1uV8aEbXxio+YyslZcY
/u0XNx74KT85y92RKsyUesloJkH02Lv10yfgEmkoGigk+Yq+4bm/+/fowssSHFjroS0qhVx2Ke/I
Cnzu/P0OeqgipdHGe+a0IhyvsHdqtzJSYveua0L418bCBoulLICsTEhL9ZJQUgL2/xbXfegoquBS
+hmQ4MWgWowAd8sLKCOxII63PAdUJe3W5IkRCXbJeK2fY95swP9hDoVArHjyXNDVKJrUu/wXbKZI
xNiOb+hYwft3FMPSvxUm0PGXW+zBbEOY5D/iir+7q0wLlcn3JGPbE0lm3fGZZ84Q+ttCkRQZn0+k
+BNJx3ywQGdHadkFdtXugz5M7ISlSd9Dd164dbpgkwk263vsfxIZPuw0MJBPN2BksJkRtxoc3Lc5
9+CGmJkdKZTLJ0soLZVfbat1wnD8p60pisCAsU7KOP3jdsfvgYDqwVF1Q6s5xcpIG1d5OYeEOQld
H5yKp1t3Skwat+XGTQ8YhB+/uSf32cjDfRFz/pcf7MUv8H2A693Q+JqK3ML6Fv2Y4ZqcMIAu0VDn
I7mf2AvT5VkZT07jEtkuSOlDYDNb6DDyLe5SwzZLgsm+tvKcBE63mohYazwTftNHoxig9H4FX6QU
KO4ecb9HG05YlcWv8qp6n5WVWiTAimWFKH0+dPkHZ9Gna4umgN7x+ACuS1MtVOy7F/TleHUgDPHC
CZ/MXC7/8A4aJCkioZzLZt4ul+LdB8kMHtSHNdLwZ8ugNnn4RNK68EEjwi5yet9qu751XwWs/n58
i4qYdqxOw/Umnrzvs1fSaskYfWN/C/plSHxRouFbTfqV1Azoco9VRjr032CkrawBI2J1tzR+S3CS
pUXltFgRtrSoSzPQUXZf1vOt1eFiCPM+jU8v0K1NWJzN/dDUpIhWwU69MsOtqrwZT+0zzdAIwVwx
o3FXgUcbZ1h2bKPONANsP6KRs7C9oU3qfqU96Zzb6x6AiQWfFAiyjEwSLBjphOfd+k0P1bfzuxLf
5HdX4eJtZ7L0w2Z87fsnOQn/wIuPGBO/EDcy13IACOpbm41bf9cg/sx3aYDh4+o21IJg6HNXZdjF
Ddv1u2x2YFhHDuWXn/9CYDG5X2iLmADveuxxa1M8M6Jx7YpTUMlWx7ve0WKlwffAG6x+bOOaNYu1
a3tepgChFYjZXAkeCfYpF1WVY4JS0Y3ymkU0YeXymEHQNeHED/ykMWuobhCFdBQNuuWux4Pk+PvW
nM2smn/l9ImbPaQM+tnZuZGO8b2fByTva8NdVPdXhV4t5CjaG+t4EWpz4SPoiJF7KIauYCZd8Z9/
/2WjIhc0ps+uiwNinN9nQPfWOQH6FcD6xOtD9eEcn3eNB1my4iigfV25DE+xN8JXyrDhXDKfgYKg
70gHcTt19QWM2qb29+1OepUnUQXq9s7p1H7Km5Fs1u1xdCijyTl6syhRTSJBXtSZIbTNR708MjQu
IXeBKMAAB2jHJ8N2Rnt3LX/KodyqknJcCtyGxh4iABy6RCRtFk51yBPiwyf6orwhLRRSWCKABRcz
Nby74OdvTchYtzBhtG+ZjgSz63PnDpzUKDtKlBdClli1WYRpJGMstUKMgKHcDibFlZqbWGXg3Z+a
zr+/W9kFZx4O5jpn6lF4H29oyWoaGYLq/pyPJ+J7ScxAGtTUkVcxql97UYKvag9UoLs+Txj1eh7J
gzW5sqxLcVzBAVWuRXdNaQtrKyO4DpBqs0T3lX7WrQYcZphbKD+R9fdPu6uTzKPt5NhSGHkDBuQ3
dEKJ7A3gTzg6OjLNLgM49xDekMAU8x4GnO32IPM1uyXLyqNibVHu6PmZczRmKSs4MrEyEnmKvUhw
YzpF0wbaKTFgUSaEKJmVftYBpeUPFkEomo9rYXTUAm3YsX/DyH9pcQlBSwttDBKSEKLlRNTxuVh9
yY3e6Onw0gDFfhZMG7LHEZZZdtiVD7qAl9Cbro/QriU/b2k4MhymyHGuLuisx0Mh8zVXs74RNOfT
J5uZ2i0WnCGa3hRgQEGIBD61Qj/tI7fcxcIfHcDdMlF86CKEnafjTfOhHgDRT4XSEHiGRiuK77p9
Bz1z+pgZFph+77dcpqzug5mvwm+6GlurdK/c5DnLLnK5zk45BQJsV4WLWZyc0Q+h9GH6oyjkOpbC
0mubbFKWxn3LlIKVdbp1C4sDTzXCzSQ3BE2b9wehA8Hj/zwJxd/JSdOTepkSY7TKpXxWs02mTaLJ
HzJMtC9OOoJ/H7y50IlPpaylyPwM1hN13CA7GfLkq3VWqe9YyrXm0aGK1BncvlS8qgfeSHlmm+LG
noazyGNIKqlBOi0FgtcQzQCJxI3BIblZKzN7gZrgxMEfTTyprUxYtu5rfYSdFjbxTGsVIJyPwsV3
+LFmFB7tkWvWYvsNOu6nwHRJDFY/MCbh+c+DMyXg6rPV7shMolJe+rH9GoI5uHdb/GvFCZbLdlkH
sbjCDPDC9awW8GqeBaU7vezu+BcY4h0LPHFBh0u9IxnCDB5Ll5CdASAPl6a67OBZLGi+Bs83OEDA
I8y2Sl9I/Cy7++MfxIAciDZVZXKBn6Gjzyg36HUtXx07Vee89dDhcHfzgUwe2XoAd1+9/Np9p8PP
zVsOazn5DkBXdH1dSwUpy7INUUZ0SBPk60g2Lsxb92B9pF0D1WjAhy5PWdjGIHgXxnO1PxkoIgHc
u5aQCRT76zX4XZ8g7WTk4Ce1wNF0kfT88w/TNJMsn/oCuuz/i+Fxl7NyFWWRMh8tuB+qsfRktmEO
H04Hb1r0tolAzbF/GhBzCgSsvqhyfmq4GqpJSIz/Aw3S+Ly7myspTzaA9p7rBDoDU8Y6Vv+CEJ+7
mxfrxBo0+sCIuf9ZynKMCvrsRUHjCcrBli1x2dX7sOPHr9pdAngnwtAd8fIHE+wudOMsNGst6ydz
Hlog3YDqke5C86yp62CZzScFUF36dSChIXeHM6puFxZgKGlRpx7gsDGiolyenwsA2aPPBAqA2frY
BkpoSX0ysBJNzW0EhxpxoQ81aq6Va3lEnNJlqWisUp4q1TqJlv5iOtProvCVd/LWPc9C7VnrsndZ
W4PEZzK2MTCBsOeBaWTL+oo4wyUkOAqrZozYislgCeWEBrqLo3K00j0SbyeFv2yZ0mej/gimrUae
K5GsD4e6k98hIvK9TYs0fyxt7coNqTwHx2RkoihBN6zpkFEC5AuOLYmdwjLmZBc+w9sjFEVMh+Wv
9Y5PACErktD67kHd0TJJQLHPY+V5Uyz3OtH7q9y4L4wPUu79NxJ64o2hrTJkWwMWwN2F8XkAWTPR
KX3hayi3ULNUQt/kqtwOp/RcO6mWAjlBOKMkg5tE0JlLAaQRLbK8xtBsDCAc12Mvv1QBvNejNACd
1KEQ/LTNc6bE5IuZT2leBLdH43r4QFaAmmwb8RI+UuLgWEnQO1zQUvTXRSgus4AJ4etMFb6jPPIB
VLKd5+GKm9TXScQaRe/TTv8T/zw0T8EdRWEhoHvvuAbCZKl1KBQZRXD0W/GLa4xFSevxU6lV3TbX
855YeQ2jVPcBs/+ioEARlU2e7FfY6Gu0HusZX5UgF1eywDw6YPKV1CgJquBTVsjClnMmW04Si4b/
LN/hkRS9+gO8AtdCBO+ar6rnFOV9JpkTK/3KywxppdyuJAOpcDzna4f5UJOs+3RF3TS4dzbBfqHk
4j4rInl25KXTCmJ8NtBUyMkpIMnPqKFXBEVbp/4WlGwu0a17t7+pyv03E8xfaF45kEtUxcqI580v
QLzKlew7wsgfXf3wtx33dBTNpaPoGs7n3OO/RhgOR/CmimwzbCrlIGnzShszykhKFhLIR1ikLCDA
pBgU0AwJ3PgDT0FQjn8US23bMREg8irDCOfE5pTkrOet4sAyf7MwNfFvLrE+aJ/BVA9ATuDFmMJl
hxVTVwxVq/SnXBG6Uci7F40y+N2/C1QD8+5gQoIf7cxETwLWVRBP16ARL2POPWSmvDgpNF3cieTd
r1u2iO8DaGrZuQK21DdGUNaFbCpWi2aXuK/68P2Ic2KEirVDBEgEWyR85Fi4Jp1oF6ymXGL1dfAG
qxY0nYuKjgAUmPFPU1KGpvvOyYC4+7GspyWGYx+39hRoR8DOOtTcY/tHpkNluZ4dcHHQhn+S7tHA
lcZ0FwlpNKfKVUyixDFK2eoRUQyy++mfU/oc+9yeFdngEOE/1TlrXli6kzWEHzoO07aYhdfCZI2F
5Q2ocVi7s5Q0KB79SI0vR1JybSJITj2fF9QmzoZGqzBUeriI2OnmBQ+lC8/yMezSDLYAEpOZVwDq
xUAW52Ko7BRPylKJamqPHTcE/qI7WnXPhwsgS4T9z2br4tXgjaxBjmgNuChTb9z155OJwR9DEJ3R
x+wmFEm6xN0W1/nNeiXkNgrU2JTgYTjiBFsI1N7B21WnkBQVSSvHZHPhaxuO7YAhbKXzyX3q85yn
o7bm0BfJb5epy4x+pvwbyxzFGi+/6aI+OTONCxxLJMdfnJT14Pm7IwchDz7oAj0/ZCkclF5zU+MS
TlVz42x0lfxK59O+fzrJ4kFwmDQ56qNwngJICqEB61K83EyWEUxT1nGrc/KuSuxfrmZ3+Nd1eaCr
EJa3Q670i6b6O0Nglgeo89Km8vWqj7dWJkinS3J2dc8Dn+riNYeB2Lhe7l2E2kcDRy0zGOTsw+Fk
OCLywRK2rLV2KCTnS5FLo1rt4kHeTip1Rd4MlB2Ndm6k70uyB6f+cpS4qadIW1zCgwc8gL5AuowT
daruSwWWQ/V8WKHV7/gVOV4Hljd6vOy0AsIKJvM8vwDp3VuRkVPWTRaWxPAXb+oLiEix1C7qtPUc
553CNySnkdbAqSRhKWlgku+rrszfCKziZCB/cK/r2LigcH+Ua7SKOW2AdYqZmfRUvWDoq7awgr0V
Z34+Yexo60uGk2r0UU73QPMQzpPdjX9cKLojcWTUylHF3ST1nt5FHEVNAXyeWUifLOx1oxJACV52
5CUpNrS5sapNSTeVisjFxqo8df/cZ+ZDasYMJ2maDNC3GF2FccRrg0mc07+6gYXYSQrljRwLwdgh
Fjp0DKnOZ+64d1RVaGrYvMrW17lMHZtAK5CNStpArASrYT9/BUbHUuNipycrD8ZPH/iMxsc9hxbt
KgZANyNN0BwG56NC2cIXyBMf8viTjcnHYpQBYQvbbffFcFZ1egaLGK9ASeVpyg/XEyE1m+eYmnvs
Oz2HSc0eA9Ab+n76K76dE1jORTFMw0InPppkr9jWLUlfWMIJKBnp2KHvBowfJxpdoahtTp0bD9zy
zTlBlR+zR++Jc8rcx6CenV+wl/PezhdbyvSBn+E9/O0eFJPG++iuxRBiYPgnxnMzkTZ1HCzSGVqc
tvKV+9cGaoKkixoaY7gcM1aR5z2TTLAk5SEGoCE65LVZ7L+NN3Ui8ZBlEAGCupGv8wJY8AW6xYZy
zuxXDBFDqX29X5hj/tHtec9e6iDrjPK2TwrpxjuUbTRvDdapTs8gqVDpAPq7nKwMxP0VzJ/nww3O
jF48tuncEJ3I0js4AALTKI6WLikExbdhLE1EyNzvpZ0ihycYmT+ZGQzRa5XiIoDdfrmpN4LTA4Ur
hxRADRafy+KkrtUeD46dFUaTtHzpCVSSjkwZKnQA4F9oQOUyJdrBU2h887kJfOtfz1ClEiLhsyn0
vQ4jg+yuXoLOfYprLZiOSCLJw84VcD42yUKSf2XGkWsz8FMIS3x52D4cozFyM0w6FztmZgQHxjPl
emUTerDU0EKOB4hE7LhDLIQu9y923o/3VyoOv/vDm7qpQeB/87tkI+rMK8LjGHTX4QABpfOfJyfb
giPsrg5KJAF3dUt5dDKtVGtHRIkqhFr7hkpCKKAFHVCgghhC46QzW1SiOqXU9TBv4LicJo1/b/AJ
RJbobSkSgQ7FjPZpsPiqLkXEbzVg0rQY+jsDwWLLQUTb7xPEpzrDzO85Dzus9ouJIOYM8BqRbLzU
UhOfU94CizgtDlu4npYdjlmQYHAW6yHtGaNgyX3cPcz5qA2pzfnQSygAd6fEDJsNWXFIiK43DteO
nSE0JUqhGH8aPGOULNLpcVCq9hGNPJ4sq/EejDreLteEi4O3YgyNmCug+eV3glOfhzIl1VjaU9Z/
o6sUsrE8EXvx82SBDFS4yCzqUXJGcaEUfGUxcfW6lyHqBeUY5uZujYDUBEgbXrxC19sqXqpd5Gyr
oIqZmxdhJGsrxdRVUw0OxSe+8XqhAO+TqeLxDrGKU7XL1qQ3u4F3wBnKuI3iyC3mJ0USHu2Jf0Tl
nes4CbywcQ6QU/WJmCo7ANvjJmsrP69tOW7iCG0AC7XIEUd8VYoIIRCSOMjiqrDv3RTqrgPlOqbC
/ZXbq09eHPQ4ibNi79hjQgPXvISt8dzZvdLR/dlfDqf7RsYWh7G+kBLc+RhylqWh9jFpZ8MikFXD
p255hZqo10qcL30zind6iAUi/oI+YbrVO5Dk9x6GHev2LyOuk/pEcbqO5Zv5Gv+CDNMWUzE7khiG
K015gLZH2MYopUNuTh2q7ovjyxASLykGrvx72/xGW4me5mLA50sEV+bxGj2yvK5Xs1M1y5T05RVW
tk0/c89FjkKQ/s5eOylefyZyGrkL4ywqzB6b9G9bVkKbJ7wSa1PIteSfCrcCobgOnbV3zBVeXSAJ
m6i3I8YO5wjfgcahbFzrpXMROpe0IPEDIEiYWDnSATCIk2ZasGxBVX1KLiTre1vA84uDRNIDnzVq
qjPUcYa2A+d3IxUvNDfHhhhBepsfn2IN++JHxfE4LNXsH2tEYYiW/lcgy3n8GZPZmqDPxkjKSDe9
OhRpCHtOaHtZ/orQaQdcFT6m63K5pIicnZ3ULtdxQB1sana8gnaIrMNxBYzSuZ9Hlany0HPSH3vf
1ao66j9sMxntyOJY4mjRfDvfYk+omkla/XwVTcwqRa2bsbKk7i6bRXG2TtE1RdIbHKHAxan3nx/B
sqtoxOoTzJ0ZXeZrk/wO8uqUiyG5MIN/sw+vvtdwgcqTQqd9Erdj/1QKgZlbxuAvBW1b1B6APMfO
nXmrlspzZ0PUO9a5rflNrF++r4/QDpa323OXGy5EQbE+8EEOZGTbQ27CsiifI8ADgHRNFW2JC43j
eNwrQF+aYjuMX/gEy9/n6hyfyx/ndaGZ1BDNbYAJjh61+23efwBEbYDCWKJ+iHjxh/EJrpLvfaAF
JJkaMLgD7j1r/qW2LdSADH/HPkP2dZOLOk0es9qRgxL9Ts8EFqh7Hz3mdqL4vPjOSA/r7lPoj5Sc
9t6R22ZxmTjziqx5m2YaRT7H2vIabTNhedx6zdORakP2VHu0LlfGIuulHI02cg0C9Eld4SREXYw2
ocJ/AetFJmgyhmqwviDBQoIi747vV73Pf9Ql3v4CPqYWjqvi+AHyelsDMyGmO7jQbCjLDuAEMhz9
/kU9i7DHENJ6MfPMSlCcMDvkgRnpQiPntGf1QnFAWNADZHOi6MtsJ2BQV55EIPBaZsUuBz4o0pmg
qc4PamYFeCA6RGtaxVDcmLFt3dBskejLV2EO1cp/ZVFtKWXDwKhkJ9T3zBkpEnA1ieYlqKJG584y
Pneqa11+4aWZvI32/sNWMOL+hunsQz30JughUyzyUFcE/pUbSQJ8F0mdcgpdUStLKUj2VUH7V/dF
oXGGPY255E++dnBL9KEWzcWECxX143SG150D0bnTHtmArYx14ITAB8BKAd/KNIP87v7coYj/C4Tp
A7fUrmC237gVmtEJnR2uc7aP+saZdXTx2FrbMBeozYslvlq2gTvDpoR7vPSPe4lVUAn1Y2wG9snj
ZpeUi8l30D9k8Ge3UeyDf1EtxeJPkluxg+Iyr1+SsRSzi/pP3QLUHo/jbAUIxSu4C722EEZt1knG
hc6DRVDjJ//hbx36arQiRtpM7oe8F+6abDZFyDrJM1WD28gS92JoOmoslevRc4qZEevLaGr2vVgk
bF532iQKohLjEbLjzk6Dwv+hGcYdAKfgxQ2UOHByZub/WIp1E0r6jzLwUAnq8zyHn6UgjrbTH+DI
2FgGCFehKcAgIS52Mw5GaoteHaXzenFNpN5aU9RQ0ZQ0uB9YZC6ANsYf8IVkJoDt0XygAifqIkXU
ZTpFU1hDAmz6nTidgAQ71y2c/NDl0Su5tV+Wb7u2Qhw/WJBAS6KGru2KCBLNpfxlxEwyw4Ujjbdd
zE3ITk7JL+QSGfnXgGVB54xkY/hVIsXrefv6DuPY3rx/6H4U1ckhQl81dn7SQZcK1zqaFlhr1rSr
nD4Qk393qJQsYcM339j0cf6lE39uAx5osL5FTQECMF4N1h1nikY9sEMvHqByzUXbdRwHMyOh5x6H
UHteIY531Wlj7dELcoBRLqF33VkhAmqszQWBsjWVbZuFFC3r34dRKq4wpaL7bzVBblEy1mkWQ+GR
FawxQZbh7ptgRipjcW0D5THVP58MwRIICn0fAmpsqdU+F/JlekR61ip3iS8MCFApcpIxft7pz6NV
zLeB7EzZP5v1DybzmImK1G3anqLLl/3vP7EksAWJJOwqi0GWp1pEXg/d6pr9NqXOgHZYfmqO2S9/
6Q5j8oaGnBknc4FJ6Xhi9mW4JA5m8hSJtqxb848unXJvOd92OjEvc96ATJHD4ceYB+ldnZATeLbv
c4EZcYTB4tRHkETljjWZMtB/clc8IpTkIBaypjPYSA1ex7XhalYmbY5JSnHvIHqqKbOqvxKVStLI
sFB5q1bvLb+XuGdhSeWJfhQvm0/wGGF0k3GPFqCv2sihoX8oShv5x8zUQKueNEOtJPIAAHA2j0rn
/+wRgpwXXhcC/9VO5eNFeQ6a/1aSNd/cRCOIAelDRDtBJgKDu53sWG9Zz9gerVoA1EMgWS/S9D7Y
lP1bbZG6kkHoU8P1s6MYBpvEe3YnDJikuT5wMwZHA8zY7YhFO3I8n9HbJgIY6YB/3yQBLoNrbLqH
rRPI3uKG8uPs/f2Y3G982oLxfgAsquhF8TgJ3nZhyc4wSPftw99Tuv4GTI3CrOrksMgaOFgjFxXq
1+xpWBWMC5YX60alHl/P3SE3awemFjCEKtVjAOh00J5gag3obRavRVGjui8KDkrQqPTE3aUddXsL
NUuIIqHMO0zCMTGKjkR4+K97Texy3VH5+yThCamSIpAGzzr7/KtzFu5K7pOA8vd0zi28gjxSgjCG
s4PYpKwV9NfnWr4SpIPF+Ccs312/g/GVY31gFT1CLYSdnavO4skbBWZpL8RTLir/ybLBgE/wxDUu
ZtRql9pNneETl+QFMs2d1MyoYWVIxgds9vauy69cDUiv9Gn0fwAOsPpsgTnFllAi4BPPxQOS/gis
LhxNMQmIvn5TyE5kIBhEdm5vXF8vVFrgGEs7BPiFZth9472xQY4qGpcPJ5uIEJY5NZMWtgkw01Rh
bnrWLLw/m45I5mXD1G/WWdF8TfYyLgIk84T4z9UJRzx3NabdMTIsLwu2rTDH1r2kAzZax7/hKmEr
h93wV6yruQbBVxCy8NODK4wjukU0IyMJgg9MoxMME20ksIq1FKS07e05tgfezysCxWVNEJjZcfO8
OlO4U5nPGcQ9I3B2nqfrarPucn4VI2I0fAHY4+kOxME1MizWdyJ0tg22x0H1/wsNMghNNIArNsAD
m4SLW2/ASkEoQaymEPTAmHcAjdoiwNhu/oTSktqqlTv4+XuEQ7xF4eAGKO/GteNKfWbDzwRnV4wt
n/vXdhQUxK9a5mfz8fSQnFo1/KjuUlZ2+yKVPEzb1aFVWVPY4KCDAROje8d0jrQ1117ck6XOGNET
dbGjRdDbynk95/rse/iQzoCylHQNM5dlpso8JZC19KT5TouP1rK0PQT4t7X55Eljf0NS69fB7cbE
VSJAngfVT6EJyTU2MCzrYSG47iaxRy8oUiDx+fT2MJZjJWRHJdtobZCMGsjajgnAs7JaoiADrFhM
Mg7F4oBl5p2gYqGcvw2dzvA6dG1X2KUB5VxDzxmYT6oH8ylcjOGWcA4H4L7soTuiKi+y7My9rG1k
VYbZGiuasjda/ke3dJEblIecQAhEZBSFYUm6FdExdcQnV0Mml7XVwr/HfIg+tsEYOFYgrB2aOOD1
FWJMTGPUW1AKyunlhrsILg8nxiEGMGMOp2+gDLVkOf114H9c+dXmg5rmpW1OtgF1uhVLH4Yksg6N
6RpJ8QzqFGzaYboNcqp5iCt94PPqkI6Rvw/Aq1sOhTqZxj7sGHt/sRauVHs56xT2whPlpDLH5Zph
O/qJRkQAZq4S6FWKvWvoPjvoM18yHTrm7tbNDoFFsH7pvXk8B5HVmHMYrAKCs7veBidCS17/JWTy
PSdYroIQaskL9HwrXZL6yeTRMuGKLDkG7BXOW42dFKTaruj4zF3pB/gb4Fky9bA+xmJnYF7eCWkB
OOoORGwbvmf9kXN8k5k90Dxdh8ESwWyJXNZtIH3dffQLsk71fbVbY2WM1PXe9dqcTzM90/ILXMFo
jdl5B48nTFBVp35Cbvq8bRBRkmfR9QKL2OjQRp7Y4H2xUKZuJOVChz0+bXHUmli0F6+N+697ZdU0
pnP8+NHbCk98iZRskzfdUgiVvpX//9xzj51DrrlpiQazAtgwXWm9QwA+rNn45bkpv+wBSQMkgu8u
alsOkCix99JwfcMPI3iuO5eRkYAmW6Ih8RnKPuVJ+ERxCBhFtKcJ5VyrzLqIlIu0JAMZSc52c9db
2nAwie6VKO91H5NdGGat2i03ztWPnEm4APveXRdKMZC0TRVyiiavS8nYjeqL3GsCUaIqpSXctG53
nNBsBf/+rhkMK+kajUsnwrIkPV1dAueY48U/vHfrLaRwNT8DBasli14yTTVH2vDFZ/mv0Tpf1n4v
R9ROu9R7H5nv8YwjkNa9mUhx3ZDH0U2IgfOm8NyNCLMMewWF66PKtoxpJ67hEhLbppi1v+cYFuBJ
oHIfLYg3ALRp11oOgYbwVPMoGc36N/DSvvBcs76YVU+oU499YizcGU4uAmp3gyyLzc+H6Az9eVz+
Fl8rmQ8Mj8CEO/bzJ5KLdUrVxfGS8t2Pae6DJA5+fEgq+5zjdBQuhIT6aBzkuB20XzAKUzM/ecBd
WH0ucbZDsFrhS+quTtot7coh9r/D2y+SA3FIAvqy1hEbiopKTq+Hjx79imt/kJk8ye9yKXUBWmTR
iK6XMVmYVBriC6UvSzgXbEB6WX3sPIlzHkIoNqFTX/ZpvG0BKZy2p++lupNu9zkBRouNYvXUqj/n
efzzt3VsFRfTKV0HVK5FfE/ZXF7haAb+DGmvfMo6MhwTTVSvbg6VkrnsLaPy0uLG1ab0XjNLakvF
ASKBaeFCAe0xbu20JgVdJkMnT4n+TxG7dq2a4/aGdVrmBXOmfrlbyQpbuNwTIKj27/6C4dNwflRb
f86QMaim4mpDQ77egtb2uM1SKV3oodt9en0dKDsrHmRcEJrFy9V4PXz5w4bAS+TmHv48eFznH2In
3udpHMpg1Jnz3Gw/rzToyqylUVCev70LZYJHturddtVh9nQdLQw79u+bkYabw9+zMiqECiy4RQ9m
qfOKWFHJmsdRnDHIgl6DiEn+QwUgMmcnYDZpH5ejzU+jDiasoAEgbr8SeCIhLQYMgOxo4L60KiD2
+6tAPuOvqvLt6zm1KFJRBEg6tIzlSOGwfuyl/0KiI9YOKskeWc1iUxD9Z5AYBuEIg/MR6zjdCT5R
XidDOvs6sxzDaU4PUFPWF2Zyz4Qen7jdZZG8IKHaXOLaYII1d6zqrtuj/IAHZt7uHmb/JqHAKQY9
9fg2vT3MuAp6IYA/ipQpW73ryohxQa447347zgevo1BqwYgW37ebpbnikFWf7OdBHMTKHQ3Y91ci
BAIdRDHo1pTnXQUQC6N3k9Zh6f+DKFo/LJ2VPdrPWN/ItqoqnpuvBnt2zly4VPLi8skN8sg+bfE2
a+AYK3R0A6fCObXWozt1soonbvxRr7NVbd/I6yIxFeE2QQjjNu2tlaw0lLAkBtu0lPfhQ3TTSrxI
V04Kt5JW9tPGDbM+NMb23ELUXrHDuYEhyZ+EI6aZpFgss+Z6R3dP+qvHNL6DIF0fV9xB4NehV8Zb
PS2EcsvJwsOrC/8e/0OlNF6r/rK2oD6dQd2M8R0rs8X3rGufhMfPcKEVNDtQIQQ0ClxEPiRyONxF
zMyV9yZYS/fBrsj9s+0sDiUU7Z+yRomRWeAo8JD5qF3gIAOZ/3uptQlxCvkbB1gbXqYlPumaoCB3
hG4HWIm81VfgPUq0h7cZvg6syo8RG1XUXqdKsDLwEMYL9/Sl9YyFlLi2UNHvO+TJ7JC7qZufyQiX
cHV9468ioSllAtsZ28Xkq2XK1XrsW3hkdDfySI5SFVv+hU3cjgsmf0qh3++dkJyrbgMujXUMCHCn
j6PWEFooGcnLtZ4+e2qXE70vURvn6spJ/39ruvm2UNSBKdLk3x6IWNDqWu//I0xgM20+AlffILuT
In3IbAu8Z7QQeJ3Ph0AH4p3ZfWOObSFQllMcwryc1szegigQ4FFPgk4Ppq+VuxfPwRucwlTM5cDU
o6/JOdT85bTW6ShD0TFQZ8nv2WRWBBx6zJywdtfpHfzrWv0YNYBr2v0Bx7ZG6aFP7YIbq/UXwVTD
PtvmNqfqGuXqzmOJxYaaq5LW6y2FNJ9/aMgpvmAaiZydAxAdazdDTUZ8Ne4zUwQ6qxenAOAWy+eH
07DctYDUfNsXa66hHbi4rnPDaOBHD/kbAlEVa7y0N6uGSoq78Png1AwvJsdKY1+uMaRkhTSR6H8i
pSv7z3vp32aH5JIXUVelTDQ7rfZ6lEFvdkyrXgO2lVxOK3uHfsoRzuGFc9ZvR0T56QfwRtbWKYUJ
YaBhW0W2pAELdyKYz5Dd90vzlA9geDTPn9X6YdbqAyzw4F4DEtIy0YDwVrITctb4+H5qjojI3fxi
uczbtJ4jWJr90jjnbHYNOp2aRgqz91ZKZ1BWraLmLbx0snqGa0RYaqHKEvyAdmY2D8eBP/gDhHEx
pniQSKODJZeLq4iHhaKKz7JNg+34M3bLKVMZGfLy+jBgn+U713O6zxUFq5oNetQpLVDLurNmBr8q
JmbHuWLYOn31NJHFS3uipABZ3QtWlVMerIi88ABhnha4HrQsneQjtPbl3Y3fPwgsxOYvrFunE8NA
goYJr7aD/tplqHh8noUlwNGX24FmwC0Pa6YxXWSUEEazpKjotWAll1n2T+Pz86hjSNq3c992pv2p
8TBEqJ4Rsq+8NhJAPXUedwXYICOqReNNblI9mYANN5plAwvb62t2lwVVtdQUP6+rI7N0AelWfhJN
LQe6Shd3lKcgqVnBNHq6s2P/Ps+oz7IQryO4naaE/0nfhBaHQUL+D4Y5jRbjDBPS+CFtN0nNKYR+
aDeBg789KJuAg0HINc7a1QzQRN3y5XoCs1HRZhr4e+R4HZ7Iltdxj8ewwnnTJ3O2tTSJP/bWyAOm
7NPqoFomWKlHKlWJGGtkJhXR0RUIo2hVn4Ldop70jJO9TuIl7f5cDj0fmMZTAOe0GBSf1ejj3qMl
uPkSF0UIC81m/6INquM4aLEih1gumNagrv94TUIQCDiKNeMkpSLKdwVOcrpaMkmKTkTnhkpQvHfx
thvJvG+FOGharuvcoJ/s4yq70VLPD3EQpKkMsUCd31TkFRwo7z7dYN0UXp28mW28854yU/HI8QKu
4y8FfP8HgDUmbeXfjfZfua9hzOzTgo3mN+aknQ0zKn9vJ8Fwkk536cMxLvG3tGdtG7eZPCyUlUsj
Xu7SYJwwIy83utciUk4tG41oXdYzMJgFoFBYldLFXinKhtGsPZlCTriKud61eZqfRK9i/EH1rnhI
/10eh0+T4joqzjnzmZ0HBp9rSQUJokbNFWq9EVO0V/MRd31qnpzPM3hTCOQJSOJ/RCSziTF+5nkX
MXopmy3MF4a/DPoRreXEY9hUfcx3wLlAz+0BzS5UTAu4CQUZQkV4So+JxExTh6ETIY11eqnsi9jJ
ciKIKnQXe5wm7RtFiaIiM50sIXapwjA6R1Osyosjhg82LhYbKMvhfVcp6mBicGOU1swFDQQcFMT2
ZDShDgZUjpoVNiaNfRgqplWkG+aWVvWGKVnh0BNWJsSFJ6FJRzWopWtZrxkiZa+KbUaGs1vmk3HC
PayDaEnJ+fib/NPLeFR+qGM8JfoSgTU0G43Q8+TfuxdOBR1MvMKDtlEwKXvu1R+OEk+6IbLuQZjP
JLSFxhQkLx8pw2XuXFetHXA1CcCXWsd/VVaojdsLmxbQbAaFElB6HKsEH55kWONWyCHQ9qCXPiUC
BN+Mb/bRm+x0FMiO3HlYxkP5WUGask4/0+RcjeJAnC4n1it6FlBPnYLPFfxfqB2ctkheQO20RSFf
Td7fZmdU5BR+GNpAxl38pYX1hGykP83ncTqAIiQ4NUBvEtoJnVXTlfumPXgmV2t/0yOHjtPFG6I0
e9UYC1WkvCuKUpiHFbAa5OProueSbBlZyLYe0giSxL2xZS9K0JIES8yN5DY+0L/XwOi7jQW54xS1
dKrA/v2NgzJVyyN9DQMZ3gtmvNeISH3PFcRVy0ez1rM7sXK6OeUnTiCKviKbC1RfgDi4YgTbFRsg
GSAhuMpY1QMzanuf44PRRV+MluPORahD4CPvmxdePYMWJqIQTV3UW68PEJ5tCUt+K1JHmnPb4Uxt
WFzG1E1r5/nxpSHbR0BAz9te1lzVTPIVVKVeWdA1IgJHg/5QVr1pO0GEw2Qxq6pl3S1NMWKqB31u
qHWdef9L7LzgAQ0A5K2igQ1CHVr7809BqXy4b40P2Zu2Hlva+QdGeEvCZRq93InoDCScE7mhx7bk
LVwQY/sNZMcWCWkbYQFZE4fLEcbzgXGcFts8/7zRpdyjeaIeOUtOOeHbl4g+CVjF8n8t0dgGVouZ
mvFv4f0Ou5efXbBIGL8niS17Jf28bxciBa9J6jVzxhanp3CruvfE5h3eKEFmuOZHkX57pCYbPivd
vOiMcdcEgap9Rdbt6fpxWZP2AYJ5Qa7PKGUgvkrHZTctrbFf/TJ9Vklo+YiLiRN2M//FTG5DAzx/
em9eGTcu2kCQN6bl6XOflhoPU6CKH5RA9rR5a0TmNe5y0eYFxZPFnVboDxyBCoYAH9AhmA48fm3G
iMPUZu0zsosbBW0m6Wg/GnMK+rVPVtYColfGjHOKBHjOeQfiLBjD8JZomcyVdOrotZkuKEpcyez1
ltnTLt3N32qMyWoUWp+d4J9CZtIfVySxM7hJAjKSu+88fGwWilN8b70D1+gyEpu2CB1mEhI2vOhp
XMCLmFEtOh3G0Bn7l/uUJXl/oAi8XdCi7riJoR98Uf9Yp3ao53I1PQKMzKbSV/c2fkSnhCEfnDL9
kd1r7kmacJki3J5P5ZDNE6+/2N32NYvSGyJytnYoODrthmIjyd2L3f4ZkuASToVW2eQEM5wv4PU7
JodEk4flZc/b1LV6n8JeU6ECVd06EofbI3UTdW3RZWXoZ+QAaU3Zaq4EyjnSzo72Pvi5rC7ixidS
lyPPOfiVIl1pBOX+r+QA5CC5pja/HSh9gFO4Ri3bXlD/rnujQD5MLb4oKcJE0JSgal4J1eptMb2G
VcIVzdcyehOF98zArZ2ZA0XkK/DVH93lwIaifwaPCA7Bs7BGGb6PMdDypOO0igPonFQxmI+/fNkG
F3on5LI03pR0tniNjJD7ylLIfF8k0enHAJVV3Q35BCeYbm/CFzrytDTJAMBaY3lx3VG53I7jkdQT
jmd0LQ3pjx1SCSRrvJ5LQ8VsTGifj5/uSJMsK9pf3tAqsKwYxIsJRgPYVdRA7aNjjF93Q41PgAaH
1mehif9EucIXMr8Jg5ySUIFK+sWm+H3mPBflvbg1Jwq4IST+CFgvO0CxzqDgkInMMAuf2nYgiwW/
IIKKti4w9mC9ApceERYHvvlPIHY1yo6GJyMRW7hS+lEAhEVjC5OY4cPABwYk2hk8405r4kEMWiYE
MArw9k/64k2brmwqW12dR7vzawe9jmejia1Lr6bC0HdSUd8wOjEjDXajcGU+djVyzzK4OqePwEq/
L9JC1syDjbo6OURz+ksc+bwe01rDkCRwyDNLRnj/a/CKLLCQ4imCcuSqZ4I8f7GSqk3ywctjiKNJ
Hagx/FW+H9v4FDGCGUa09L1s0cMqyUIeWBmBBXrC+Z570suWOYIKk3nzetHpxtfh76LFlDWE7Atr
SPDbCfr0vbvQra5hR4I5u07ynes7EZMks2RN0k31cgJqVehLQbb3qTBQi0KJ/FKZfRRktjM6hu1R
pb3bi5kgVxohYkAjs4ipICxyY8Y4bfRtQhf/lVapz5e2pc2EkFs7nbGGkj+JMQs8HdvQSDSr1y9C
iqct7PewoMy1r3bGEUVur8qMC1TW5QyCJmHsABQzhk1tqy6XpLS0O0VdYTQ5q2SN1T2g/PUsPOA4
b8QSNnyceu/FTJBKtVR3Z2VCPCE3mLwAJoCfSYBL2fT0PByRG0G1g9mWj742aoo8Pyi6wRknJ5UN
0heAz5DgbRoZ2SBhY5r/IRMitom1ynxONKRhuEfKSRnwmV6btkJ7hTF3PlcLR5bOiDPg0a2iWm1S
P0doiKBdP8vuObp6xkKMntNowSrQ1a6Apu9iT2uk/KetJQ1Cp93ls0rN0QfvVrFONFTK8ZhC+xJe
rm+fvykzqu1CG0Bi+QJHjQ42Cx2Sw9hX51ysID49YlonDp3u86Pnbh1NSPMwgmBJsolEin17CUa5
Mp2HwHgBglxmakCVwF/aL3EoYY3CRf6QU/TN4c9FpyrZWk/rDdl1moqgraYhDymSOePIw4tqP/zq
S5abm6w2HFFSLVsiEcrvj+YPLW7044CGAjJ+dKMZRaux+/PASWJFnQUFze4reY5GkPQsKIMJusEe
/2126efSyhJZWuD7XWDd4diJu5qOFU9Asf0mSO72bmwGRTOCZ3DMSTSAc+rR3BrUVANWpjN0D2KA
WeQrdLTD3NxmwjuA182EQn8CVQEIbzfxMZgI6XUiJu/uFnWVC32MP94Gnt7hcCy5Yx1/4BmrdRFu
kFUT9s4ILETC6nK1spNhsag9UGFD15UsB++b31qqsX/BAcfjkMv1I4MJnWHwSRDCp/ame+PY7jO0
N8wmHQpJlRzp68boxdD7e7UyCvsJvOWMJowdgJQciWsp2A3tTR9d9RV0VRhq/QROwPfr8S+7F2XA
205N8qJNVXc6xKkPSNT70KzA6R/H4wbxmXJwHTyYORsHgR9+3rKwHqJMRTkWCrmQKOUpehi/Q5pm
dStc0Ub7iSB9iKi7s/9BkCHNSGDNrksjhqGkUXlyxEsy4JqC1J5A2smGK19F0wl8mX5W8VcZN6wm
/XCegCu9gnd5LweWhU9HXNYnxd2rxV4k+1rtgjBv8lJDxqdfO7uuOjBaEayUjvrQFhJbc07i88+W
OvMKrUJXujuV/TnF8n+CBmqK8bOAft7ShXB9qJB1KxXFk5Cuto85j3FqwripiBn5SNPB/UdiY+Rj
eXlHZZuy8TIIN4KiFsdNBPkUydloXYo04JOToSnmUfsr7VS1Zqt/TOMQS3onTyjiNa+sq3AyQjoz
Lt/OR6uOrjrYMyrAcLg2GA7aLd7e2mPbAnaYmf3ZhmrlkN+zZdpRdOHJ3A0MxjEillTb8CSp3W7f
g6i+DJIlJRCcu6eHRt/4WAWw5W4UuNagnIw66PducGehsCbapSkNc3Vq1kwDLSBbkYO5Y8U0PQ2a
5diwSFQURfLghDk/XF4pLa0fA4rnaAfO8P6LyN5Qcuz2xhZbbSlEIzRSyU8dtVix0w2r+XUnSh2I
JKOsczSl2hGnC/E49Jz5AfM+Eb4MEnFeA4wahxkgbi1ua5du9cwACtWXr+u9MXJJ4T3L5vd6DUfE
qd95gC1xXFsHR/oKUjlgi44eu1tCEWl6PicF7dI/BTt8Li+ewV1ygLInX1R2IcVswGcY6MxpQ3mQ
327MeyenMJ2dqg+ZFyDtSBgiga0HZpdx/58D/qWXJTcc4UYZ7s4xQwFqQqLnUpkW+xZkIp6mlxFW
1TXd1Mg1VUt/GGeu4FYN0iLhg2xgiXVkEWS7K/pFdJ+HtzKQzy7p7J2to41PWAdy2B2zT2uYAwGa
Pa3CAYZNa6GefB89RxXGxcElRD/3NNkx2phqtKoNVX0iSnCVsbR8clKmRze62oS33LJ5SvAK2nc2
BX11EDbH56Q//BBvAu30GIpDMFkN7npycu2cRGeFnqP8VX64TCryaWFgA5huY9e2JHVyN1tc+cSc
Nttt3YZxKKpFwcrfb2rnTi3UNsb+vusG4DUux+ibTUlAAWNPHRSOnwvHjDxoKx9pwWYU/4j7MNOm
NXwtfa79O+wfrtmEkN89dUZNnrzmq10ah7TUqLXe53rtntcyqOaI+WLHA3JFqUN9xNUPVWeKFf2n
L9STylN6sNWSsk4Fx481azKry5zce4xRW+GHIl9qBCF5oPU/WeeN9QIxKCLOx+YUwH9rwDz3XfjB
1VJIaMatZVtP9VSVkZw/YcTHPlzWxuYu9fayu+zhCO/gseLdDXIeoBUnaEReR+THceBuipVBZfHD
kH3L7sUv9otDAAjuHs2UwGD1N/dI5PWLLBiH3EDuKbT5KdmuWNbzgaFGN7nZ+/Od3uOINZkyLcgy
KAR3HzlQGsvIdVQohvFFd75pSV1nHa2K5KvXJkwhVK4VZZkuQ76DMY4OG+c5gYF9mePo/KW8mrRX
FqSvvBkiYEEFG4TW2/2sqlTxpVG1RH46+adJt2MsPZSbi0a33lN3Qpwfauqo5RnE6cOEuM6f4yFZ
6gxuJKSF4r3dw9saLLji8Q8BTFN8gNcf9R4qXeAnUVN44c4FVrBZA5rAQy1OkWYyBXjCu0blC6Ee
gHE+u3DwBM1nmJZrgxEsbjiRGZ/N/FU0oA2M/7wb/kCpI0JObNRLhPPcZJW3IdTAukAvrIA1KW5f
YJ+Xu0U0Ssl22U9xsjLvK6wVyIBhoNsVhiqzNeO11hnGCY7zc2xBQOojVEuaRYbJVzZ8uwC9WzlG
/Ls4TqCEnkZEy57tmKv7hoZNc+mRjY4qYIU4q0haJeo1daz5oqlVSx/Kn6vPwfn5r+OzOsrzhjf+
HwW0YW3NhTVvJvLDxHtvhWdpWvs8cuWi7th6KIDZtwOUgfHIjBJNvGYZmrDGuaG3d/yjR7bnf5Gw
03jy3Iginw6UIR4ocTO1M3xl0ZBC0XU0HBegbXyqsuqSXDE8aa2LSyV0TLV1+eKkHdojt76O5/v2
upeYy/u0bja2RB7AZ9OXTxBqwH/0JQxoa8+OiyipDsjOWjGQdwd+785BBNZVvqkkJy82Li0R+Fib
6hmAVWrO6ph6Vg0MlcnWopvMZCNwvA7zK64s6RiXvlnPp4pxC34frAAJuGF2gewokyzZmAHx00bk
Uz9X2jgX4+Pw12evgqHJRydxL3/zfQsAkHt9yiMHkzRVvON3WB7qyMC2gZ5xyYt+cbsHaMxi4VhP
tN+eij+BK4EyauoCftBdYCID8+ClqQsuBjcgMAdSCb/okWUPGkwUix5xaMyDkdtvDihz0oR7wqfg
4pdH4vkzFwyWrlXtic0auiHkKelgLhPI2Ojak95JKyHiK4gvr3dERxzDQJ3brHQqh7OzR1+/sPTO
PUrMRu85oKqC1miM2kIjioh8BIGNIzxzmIqstrIyU9+qYFL2JB1Kz0QOnMg0PB2GOnQU+RgLGC3K
rzbE6bVtPngYcknGwifL5Mk1Jdyb5I/ZvBkRWFo6XxVFk2oyli/ukljQ7tly7SzAKmJhJwHRnMw5
zuuTuVVSXmsDpWW7o8eNY02jn7yS3nO45tJTtEFh1rWP2hwiAf6I6gT+YDmE9vjG2HwZ9ppzxaeW
JvNY7I79aawHZ04Q3p7btYTQmQwgJwVfGTa+Md/BbEe+cfEgL6KnXwzO8i3aL3HxEiy7Xe5gvuL2
kxPqU1mTU2QthonCojv5AaD4jj4py2l0bnB0FxjZ2MK2ZFDqyibOmiqwrdkqG+Gq4s7DGmpgI0gl
1ePjiiDucfdZSZs+tQIlKfv1xZiEySjesDsA4+5wCyYMzYaZj3v7V4BXu1/4UIJl3DvEHrDfLs1M
ussdwJn4MZjohqdixP4Msv9xhVEkRTdCTC7ik7KJUz3HWKPoWuCK6lf8Hi3ZQ0RStHf8BXB6BMKF
HIpJ6MoOrYfYnK3WRhMo6yktPonQpzNpdGocsRL+MHQbTMOOCWdyzVvjClce4ANANfoym9nbiNZg
b9g60rXz/Ywe/ZZAWWbeRJHcmqK+9cQFSlSpKJcX7CnIqf5c5J+29VHyUBQK2boDOAV22hJ/XeD4
eTev0+Hug0G3wSCSglmmDY1q2GiqOvI3mgXHfvGC4t6N1PPbhG6jx2t6z5PeAgbrruhEvDm/AoZU
6LQPy6oEDS1xB1jASzmOEZ55jabNtFYDpbDV/AkiJ1BSGpBhnWV0dSv7xHqcD8FXM2TB557dONL+
+BLOWp14M6+QEMT1ZGbw5Z+aeALP2lJtL889d6cDDwjpj3We3rTPLLJYZHcJf4QUksz1NUzqW/XN
C3go+L2dkiVgS+j74x3nXzXCFWU97fjEQ4xVkuIz2IejeoOrP5SIc3fE1yHfI/z/rgx2mnRKxBZW
sE9FDHl88e/Ix/lCZwr6ifHRl8YMcjqNy5g0D8MyISaQEx3gQZWwjX+5ocJjyQhnLlm3CijcDMwx
R1ogku8O2TgifzY+UaDYmOFu1UvGOwBOmjD0G1mIUqJcHjTRxJ+ZnCDvjFYgM2P201Bp77yp+Vj+
7eRj65tSPJo49jZ8Uz/TIqJ2uxiBx/ufu699dLGnrTYA/8B4jZs47AxZ8OlS9ftvkpa5KDgtz8Vq
kI4I/RMy9Jfqqhae/gTnftY4ruWtVZsbfYwjKR4RJkkKOyn58pHz/35026PtkpiegZtmeln5kYX/
q8+/FHh7gc6uU7eV1MeEPRcSPb75/ADbR8gzNGWCU/2fgyypfgRDy9+ZSVHb0/m3VQdE842xE2og
gide+jKeaAIrpb0BzXd+30T3uZowdugid1bfg6do+jKDqxgbxbmL1BwG8kSgngL68D2RLE5GmXCr
kR6GBNauwyHtm0BnGl1Ww9TT8uWyL66rpwosgwxDgRD34+a65ruJWS0zDegLi1x8wLkT706DMIHl
1CaZ0fk2tsroTAPW99bTLQv54g9olfBR/X+qfrVaYA170jHH4efpWwQ9KQ/hC/ojnZjBacknBVDN
7yLLN4zLOmdqiTmDqjdJ5SOE5Mr/2DRB9+zQ1SNPp4AH1AwbPCt1eSM/b9Yw/VZqx3EHYAfsNxJ9
hh5q4skj2UbqUTexQATx7nBkWVwTzE1zYyZupxxlP5I+8/ZKRURRr7vMLAnoNUevbd3jm2bxHDK0
baKDpG9JOMfaD49fCxT8DX1Ylh/rKww8lHo4telh4lNdcudHsSH1Np/TSq63GzwNKYyuexbvFXGZ
SNfzLfvl26qANI2b6yW/12z2DcqJDVit4eVGi+Acr0rACg0ReIJASSqIL8+q7RDlr5C9J9ONA6id
2IYnxN44xHS1ejOI5YTRPj9uSkbIVbeqdCIWKoNfDz/I/wNNHGEZtkkvRcO75qU0EuTwaCVxrS1L
d1oa2SzG7bhen+Ax/vqXJpA0DdRKVR+r8J4g7ymrDsUeL1kg53uqmowz8/48NmEz6Aod9g0IYvhw
8r0H7pr77dPeLu8tQpx9caXvVQhS3vQRNf3WBbKkqwSzgicv02sSf4RvryGiriBJFExRkqFlZ7XW
lM58wPPLmJKxS2kAghDXm8t07qg9d4K/fXC7Cn3CgydG7ElBmWEjr+Ar5uMSgNe9v2eHtWqIKMBB
A4/8vhky+IyY1QeYSSqGHAPkHeN2qxWZQXCRNSjJWg1pSQfmFnl7tlNAGqlfASXahUMRy8SLlvFn
q6m7sGZuWNTeP/CdijnjuejQjX6YPuIkIq14J3RD0ZlmqcoQwL5V0FzutjoOxsfyhyuz9CC2rzRk
kczkUvrXeKsMXtrVIZjDDjfk7bldbDFidvvXPCzKn5MJfXUuPuR8OkVkJ5dvY2JshT5WpolSCCoR
NyrkhX/i1jzz/GmXPkfHKv2RoLTvV5Y3qQr6Np0iNy6Zu3WZ1fSku/ikuU+gLuUmPeL07Th2a1Tb
8ZM2XVlmyPqIdRC2JFSZL5ajCtehhBhqZ3mVjGbc2xLZ9QM3/VrjO0o9IDT3wJ/B3SBy2yqS96SF
qIggwaXwrgLDBhZKowy9Kr7c+78SmkquibgLUx5vyU994DkUObRB9PYc/KiSm4g/dJh0rElDYCCq
Kzaz0/kn8/6aD/WV27dTlf9NMlAR/7/+FIUEyASCFivnxqCCiCCMTHFUsbRxbbwsJ24jNrWU/hbp
bn2QFmxqDmrrirbRNc9R3dFIZs/C+iSm9hCqM/kL83yKyA4DTFqjunleB2ZyL/UNHHq/KKoOzPJm
GHA8rpAYATwqGxBQ1IiBLsSpfcKPfQzwoyyuI/ummFW/nq4i7uYA993vqQEXwzmTENCQxDX43JIv
pRvm9S0+697KZ9k5gSD/skK2wlre6C/Ouegvfxq2WsAAjrbVCJCNluRgwDboXshMB+6ogfs55NE7
eTyOLnS5oAfrUtbjUZptVxi+rW7yBISpGC5g58DMWDpw0FGQ2q3MSvjOdMSeZGDws6c0ulxasNQf
uIemUN4W1JmXCsgcmmMZIdUTVMrpaJUnY65zEpP9CyiDWZN1mmWC2Yd7NIUgZjg+7WvR+xMyR7kK
lNIxP9tBy5OtmdDjMfULGs5AToiHqnfvdAfs5+8HdZR4CCRHJVcM+ub2zv7o+vvz3uDRZ5qxUSyF
VWuUH/KWN1dztPAOljDAWlL3IB0g1q9nPafZY/CpwNSOYJ5V3p6Eg76ZcMTCn2CTMbB6Du37jNSn
UH+iYzQ/OSQ97PlXvU3kUd+8GZg0hPsEHgTj1k+O5OFLyPVz+CVthS7/c5f+h0hZYYE8QpQL5pcc
WeRcbj6ozFttTgYiqzeImF6DMw5NGOEqR8GFPmVENlxouWic0yiLA8DakA7TqfDFu7fZigloCIM6
SGaUVIWFYs98L1r3V9PX64k6rncTN/qKd4jfWC3RFUmlff002fESqz5QOA+Q+9k9SXWab+o3cQ/M
oj2CPvriPHy2I+5m5bB/OxeIBmQ4nJgB/zs4YxCUFKIJI0n5aCwm+yceCjWvBMQ1sFGPKSmkNjZR
OSZQU5UM47j8bQk+2ErYifnZhSXJR69Mr5mX2U4wyiay/+HPXnGintuAdvp2NZ8+dSaeYAY1Gvox
jrnYQKdE2fUU1V7ugktLkAkkGecEOMon8ghIZwI8rVpX8HHqojAhY698J7u9HK3ZAMVQt8cp4HxG
YnaLqmVJnDqbUlv1OjzuZNfK5UnqzI0k/j7htsN8PZ5QBl9nlsfgYHnjN9TMtC6u8HjSzLu54AFN
KsafxKHBTT35XVjyVcQPNXxB/uB70d0pCW9lLfMkDv5VMmYaW3MP9lDtk2qRwFPjPsyYekF1BYOh
YRZOTtqZf7co/70NTI/oi2e4aMDD3pNYRp5DPmheNxJgz4ZNqBvNcPHUZDxW6dCElM/f+DXhIkJu
meXXLk0k6kWV2bZadj8olk/D0HaZylwti+4T7oXV/0O9nL6OBi0qf4imqUNiUagb+GFEt9FBoCtj
qMi4FyPmwgCAr9DYhghazunZkdbYFzdvYfRCcTUGcEwcD3XJ1P29DZYZwB7RZauXFmPCfGv4S4ro
yuC1nG+81C2pM9V/l9Qm8jxMnMonuycpsf8zG+HRAHlfHIn0KNddEkpkKoRFvaEax0jEeVKyHmi6
3OHVVupF8wR5WHlc6EDFqpjgYQMRG9kELlqbluwVtF7vPdObNLonHGaRd30lEQAtlGd37n9EcpVk
VpKtOqMix73PT4FYFTcPQS79z+itxNV80bN6Vss83tBUQP5EcPdMKUltw6ke0365CQxMJOaj8MP/
SSRR4WV9ZYsjJDC1i2lDT6c37/fjt9uBB39/zKsSnKaWUj56PoGXmsXnPL91QEpYfk/hCZ/pleHz
DMJewHykCiMmyyooWXOLSTbNrq0Z8GVj10cx0D9jrCQImRXnDZ37r+ut1ott7X0aNJpfToL2M2Zo
sWcpJTZAWjfUOpoTvKOVigD2xye3K8oeBhMoIO0JpSjlmjP9M2mD0sIVdgC0MtIzMYG4fiIWbupE
a4xYyupbsxgebAbnarCFokiMBVAa6K6/vbbj48wQE5wPzIkXfA/0XLebTh6i3xADdGM2WihvN+5m
tsq4rZ0WPV6T7ErhdBArTY1bc5SNcSvZaUuv1UTuhQCxXCSwlxfUYBQfkD406KcdqzS57U5k5G7F
Yh+KiDPnf5H7WxuOYpX+tkVZPrzpHsZU8Zy2jCkxJmbcP4RQzUXr/85NQYXvj7cegw30DkglM14L
pHgToY0HLJefUXQ478nKRRoPFfc+iO1pzq86IFuOWrLQT37YTZKQIzR0NpVbr3CX9AQmsxT7Zlgc
aM+gj71yAcw3fEhhaClZjr280YC2ASSLFxNarKRda0b/tUTXNc5T2LSqfEHX62AhoQ6gvDJHwbAe
oF5JJLK9cCQ9qGSUfy0H9P9sMFYp5cFBp9ZvsgRfQFvwJi+46GVf7PDE+nurNuEJXH6CPIfuc12S
redqkke5XHBegJj4Kf3d0DaBZwU0Ggj/M83UBVvruXO2q+/H3hLwrHRkahqQ++hIX9SHGdz13K/8
flzcNP8QCVur8UxEUCQ4UAoeZyPD1mPyTyKOnNY5e5dE49mShbjzwwVj3YWKaG8fdaGp1/34COWI
Stbezn2d54bRbx/TAm9syhujzivxhj2GKOXY0aqpT/HajbWJsP8eEn9KdMNjyKeknsdfzycsd/XR
wsEabvZGHLIML2KiW7FQ55aRFDNux6LQK64f9sAFYjhZ0T5hHlC0tKh3TzuJsU9BIL5ykk3OEecJ
xP/nI0pgRhzITR9gOVaJAXI7EUojaVP+Gmr2mtSL1XNAP7Nx3FIK4Z1IIy1JbqYGJSdLnfvAJyTs
2HrEw0xmn6w2DSxeLADB7ag9Eb1eaBB5wXqoF/Ha6XJbJOL/SFkI1DKtcuOorzG54wCenNcw9Rno
VvNt1LNHqH+TQOfbeP9eopb72nz96FwjUUnL5aXMT2jc6oPuxdhx2/uy9E0UbauT64D2U6d584E8
SqFxS4dAZwejdp5YY7cAV0akjZhP7Msw+uLf1YLQMRxP1s6uRq9mSd6EyMCd3ZbKidpP36zDCuPs
3zuLE/YwOTFCUt1i7jo1/hlb9hg617THGHzonXsbTqfNhsFgrlMvolAk3JpeNgNQYkw5Z/A/rVi+
YAO2W8qRv32HMWbvSyVDNKp6x6/nf6hLapztT4h4uz1rcvuqZd3f67WxkGSyBbq+PtKH0j5E1zpG
aWppR0ydxkC2WOPAGKJx5ES3wiimkKwYI7UqKLvKdE6Ky3Bh84iBuEJfdfysPu9U/jx1XMJJYBuF
MgSUVt/cEzQDXE9NrO9y5B1GTrRGrDCUmTZQsWetq39sSCNfaMrQ96u3sMSXSV1oWmTRWbC0XWhI
nOZiUsb5JyTewyQ9wt0vCe21uFwQJRB5ikfRIs+8MKpfwVy9Af/vciceOodBOZMUHbZg5rxd8Hvr
anf23hU8QoNHvmTzS8kDWE8ZhdP9WPPfFmoidNJcLvbxsrHXeJn90fLS+qx8YH96PJXt/2AX3+ob
mlJIGHwDkYPdZ7Jw/oe0JZlS8KOVQ0SQvOtOFEX9Werra4JWJwEuXIznmNK84HFHc78BepZQqGDO
fnUIzA7sueSlbiFfWblAZyntlN61UzgE+geztAzDRshfr1onQDrTmv2QnJa94TNxZaCityMHrokl
JMLlHrA/8x7WWLX9rjUvQ+TwOxA62szcP3Z2gU5H7dgfJJ1h3CkCSYdXp5YY/EyRXpf3xElJH03l
pavTvYBoGUVSSrr8TwY7iTdxSYmXboN6xhI2UXQAdgZuMl0RC+3Kdm0+yBKr9x24m7CJ+YkrnHH7
qcF37UZrErl9iCfpIfZTyjNwzPdefKQpAsXPfy6SOdJTowhAcHLIMeqvfzuMYiGCEq2Aj3BB1RRZ
knqhkgDpfavRPqh50zJLawrQZ9befJqUsUmPQ/tEBZFQRhO13J2A1NYbxkQbc3kjKDjZmMIHcQvl
CAm4/PCZLwQvBR7h6EG1keLKWvAuty24uZHobiYOaXoNap/Oq+dtaBDVtNRS5gyN5HHgNNiV5dum
n/eDuPmYTa6J1UCXFW4zTPmipClchyccrLMXpe4F7TY6DDpctAKIzigN0uXVDdrNVcUafekP3Otk
QsdoUpxkFbDYeArZ670CiJ9xXQqFkOC/Pua675ExwKLfrhdzsXx6Ip59+dwZcstfwUUjYSgll0ye
DQyNP8JAtdWTLuZ72oxZFsqsWiTB878jsDy2UdUQFwXNFWXeA8vV3t+lnPvBJ0oCxRgt4rBb3ysO
xjd89G0JYQLP402fmzK9VHDFZejsWnH/TsXvydpIMLsVVeDq4J7oOde/VzYfEGReocGRsu3nX55H
apiCwFFNNkEg1W3VZKcUsu6cPU4x0fqfBkWXZWumkz94PSPvsMMlyBLV7buwc+jBX//rQOf490Wh
IgZmfbIof/vJGVt7ywkiflUxYIbYcrt3Em7eF4434RKBDxPDkDqRsUUEjp7z6OBQNChbJstJwHcM
ipk3SMZrMj7z4hrYEVC0Q2CfebJ2SDu8ETLTrDS1DBsv3xdmZ3+yKO22MAvsA5jprGIdR8WiNS5q
0Jagzsp5/G9IYOzC7KSt3EZk5oYfCkgNVfHU3pS2WE9A8etLfrKUr/VK5RCrqrZhQex5tFqTx5Qy
UT3Rv5Equhh9IsqYc9uhl5xcpAro3oOvTeFeKelTv5NWPWfrUVD8Iq589B117/8ZCAAu/FIR1msE
Rt9ijUl43Nxj+swlIu+ag4skvhfYivl8VP6Glm8Kf7qLqNrOtkzPBgCcUyzgSBWsscyAV5vJdMAU
j/R5Ey+wbWpUKZBI1fEWxU3Uzo0Ju/RWMhCwbfjS/VjjCrjPcO0Kpkup7SdFvyoToNJ8kpBzbWg7
pWp/7oLQ8m7Iv6HcOeT2lIZoaCzT91Ft8GacVEzLzC2PjstKFlooXtQk8NN0+4mSojZrbKbMexuh
N7hWi2tM5dhUgQEuqzNY9I4H+Wi7cOtqz8YQvzunATN2V9Z/4bz4COl18qZzFCs9E2xcw2TNbQyF
3siM1mrhpWG2OM9CUmcwcYUufSVOWB6zMGvSDTwZrE4Rfx88dgzuiQNSwA9dPSghZQJyqfe1fSEv
TFJarR3n6HB4wCI/X+10GpIta9RBJkBsAXn1Nx52Hht6JtrxXNxDeJrIXDD9g7woCN3WWyFSgsDp
zJ0BbKwWg1oAXWB4yWtrbGwlNgHnwi8cU95F9XkdRCpOzB2M/TDavaSl7YGJ17a66k3Jd0QTP8o9
XuFVBbg1e/UFAk0sqUeNgt8sHd8iQQzHedpeGjysgfLlXlnzyKPg2mRg1KAu8er4HPCNXcVAYDQZ
g9fpPGZUf2U5c3cgCyeJXkoP/UvL2pfyHgDRBIMCAz90NMEvxZl2pgZknAmzuDAlRck8ZrhWMKIw
rV284lHf1O6aAu8xEf6AnUQWFTDXWH6M+5YQVB/lCFdUAv43zcmzkakFHBMfA5xPHD94J2HRjI2C
50rxXbiscgQukFkUqdVoQrnmZOJ4bmlonY84r6MdlXJ0XvfKR8NoYvVqA+uHNnZNJseJHJ2rMCep
oflbDp60MsnFL69E1Sje1YGe+HfNjaH9sSPwURwXojvOmWmWmQC5RznjVQTdFG54nu6n6OPqnHxP
ohesFlQQjju9PTiu4Hr98MrPxC+3cYqPoehzJ5rZEs7R6J9m5b3j1UgaTPxR5OlxXYfd8RyPaEZy
QBZFTCXEQ93fCy21ytcHtEHOP7l9/YGqFYZDxB3d5vT6yIYAhuVhUDHFL0Sp5wN/3o6pWQYmT/M2
Ud3SNBH85QRbmPTIu/H5VaUGHqVk2cbJutGaivErL/3tgyPKEY12LO85omfa5NSTLL3esEOfa2th
UZiykAmkXl4UmLLl4gwkejjnBPsjnYasSxP4/7krFctkbjhVHvfsMWsmiQIEC2MiqoudU/Wnj8xv
GBrcGC8XgHXlknwcoWOsWHc6UR+EXT4IfHfb0WrTo+12xtgPeJtQoXBuD6hBv7nq94jnYuL2wd5q
ox1koYu03Xt8ZHfuxje7B2ycm+6YMj0OedZvxEryxEte723gjI+9QouoCdMR+sON/rmfnWEH1QHk
F6PvtOcDIGt1zaNs1gJvZ+D8QqeYUeYeZnezNSzgGBHuCZCfk6A1we2H1dfJShaTj0tnw99Jseli
wg5uO6Hux/UE0C6PkWfAThy2tPN2r3KTczYp/SZtB1wLeu29ZF4VKkRgl6xH3ALEdM67FrkfxZnQ
l/p94ZcJXrQx70KeSUN1HtU9PxkBNfI+85AfT16S/3ekUyC6iGrdDleBdSBkoLEmZwOm2utY+TSn
64UYY/boWd8Pe8N6S+cvjX7KyPg3nJBSFSOyAMSomEZ7peBBZLE6ewiY6GQp6+EFnYjwbaEV1zEt
qO/Y5ocPekZA58Gt0Ve1/ksZS70D6nLLZldJU3bXk+F6iz+OQL7Ue7QTIC+GEnA6Ck0ockr7Y/zY
xu884+uoNmlNIOT7nV3Ol9RMrfffdXtesWTar/Htii/D7h5B+oSED3i2D1SsH0t6oo+sOlG1Baxy
FgtGkqoLwkSZTtxI0Mxt/kqd6j8FS17dj6In7Sf229GVRFU1gUfVbErJ2azg5sUB965POfTiwzDh
42EzhPYMJUd6ZbFYf+1jGUXtMwoYiM0iA/qCW5mP+0dL8sdeIUyTd6mCPXHUxyYTBuphkv2wtIsI
R+XUDj4lXnrciHc4mqQ5kw665IH4oc3noc0gituu9i/je9A5+i73J0sT7kkTqkr85KvVSwmByx7M
rqevVZ1vxVSE0NJIDJMU2XwiAzAfI0xCXSJQfaa3w2x2NqOPoQCQDKNa4kdlVnL4lZKzGgxtmGN3
S12NOGmGwJM9DuBVrCcY1TPD5uTeN4YMrTc616M1NI4fcNsMJ6RUS4PiyRJS0qG6jsBpTyuZb9Q3
ssQ1doxCogvUmjkixBueaxWSN6my+3bxB2Q0VvVAM9YtWybBey3HCuN4UNaXZH+YXcypCUvpnqVv
ww/9UsBforpT3NOEVQVCl9Zt63RJM9h4EXd4hpORaepkdA+lYLHQ4iLRGmuYPjPLSgUTdAwRlnAN
xT61iy3Br+2XqxEjiHIPU0w7Oyue8M1AKm/nly1AdNXMOWdGOdlvw5jb4zjFmKMpsUO3DggOZbDh
ljS5tooZB0ZmpTMVt9xI+37V0Jzs1y+IfwlRXw70FntA/f8tkSoBEkiIWtR5bKfYRdW9uC2P7m4b
zKGXcU/skmC7XKg8Gz+omNZNglZ9w8vzMR+hVKtoG6gfZqxs6kGsDCWKQoQzmZbZASODghhHxvkj
lrBnmWoTi8n/45s5NWISVj3CW7teJM5EUxsAkn67Bfh3PwAyHdyXLuTGxcFicwptBJLJik0r0CJt
3rf2SG9p8eAuS1aQIKcA4FRjSQYP1FdOsJ8CBd9TmV9anR7HOne6DvXC2ADA/6dSvOgQ3kzcFxO5
waCSqUpoIlvzj9BbPDGfW31ZTWnh05daBVQmYKUgVyLBcHGnhX01L8d5TanFk9eBC8t5PaEqA1zk
1Ak6SnXqOCZdwMbJALpVENV7z5Zy7TcZnxNQUI8widHn9wPldCdQ1jzUioc1vhf9IPmrLbKwbS1W
IwgZEf++Ck/LUh95ecbWxQpBGuR5Xb9jRR5UVBDQFzB8psrUFW2QUPxf9Y9F4JHkiJLCwx3OivCW
TIDB3+kxSvTewGRZ6JOYT7ZrbI6+pVokOMs3KSCRqYtWLh5Z4H75ydFk92bmpEwek+Pkn/RU+WiB
PI1iVixF+aTg+q9X+Kuf51a/Xkivsve3efoA6bHulaz8hyjz2hUQHwGM1Pi4OBo0pEytPAmUaU3h
Dv/BPZZWWnhf46tCbuMPP2jBPT30jw+0lhmKGAohyTMm2GiFKXC8Bzqz+VCCTsE7t103xNGD98vQ
pWqZAr3EIpQOV3vDj/mVXSzTNYYHoTrUKnNNkTL3dasRnOAahLbKQMoLFuxqHq9txJoz7K4toZVF
7C8W3RVyg+pNfmH/EBEkpK3UnyFyFWyXu+T9PsQEiunNyjLlplqb955mN8EX0OA246UPgz/KGd83
Jh+RjOIx2IuuzqzlbjXNKLnu/xGRGOniQw3pe/7mHP5IxMWbWVuUzoxE16aikdmuh9F2ve31U8oQ
eQ982nLIfXqvwg4+LfvpB+RQCzvVIAuz7559ePllGh2Mve4bB0x2WEGVSpwxw28Xau0DnXjwM/GQ
faiYIMYoxwFL0QgSKYz65nb8qTzP8NsYT1nd6twIMBPlBuiD5j73eo1WkYGq2ipsYixLz/RVjR1f
sPuWTSNt2G3Phl0nuI3SKYi9NhF80sfPZzt/IBCxwOx08t3dk9BvapoK9mlG5IlsuakyNB+qLATZ
OZVT0roxiVd5GAI9N78sOYuqrZAjfCmLpCEMqVVDb3HXcWwfLRW7zg8/FNde3jLyJAWpcL0l+ka3
cAY5E3H5Qj6I8RJqf7S2ro6jYwM/kph8/HBMEsd8YNG9jakokixV1YPqKspvDzwxbpeu/VQWylmz
0thuJCWEjoJDLnwllE1flM733peKdPO9YSFcwBaduY+nu80XmQxFgVykXyabs00J2kSpGtR9ymPe
o6YmvVJO9PzR1Crvq/JD0frr7Z9rSm8BpAS9oPiw1iLmaNJQnTE3der1gB4n+2aBK7hptWFxd2Ge
KkwQTVyYWlr21saDa0ThtsVC/3Y5xWw9b+k5pCKzquDGc8+FwTqR4aq74HVN+Ua6ppB57UIjKjPc
kh1LN7Jy/QJJnx65nliJXxIZH7gbQ7yt25wolsUGwU2nciXqlUJb1zN73b2pxW3oAd10c/HzMvoD
8wj6DVEXYyEP3gWF/vZtZPJR8l0j3RByPJZRFpGSb3RvKs6Ayb+WCmTMrM2CdK39nPJ+0fqCBz0W
mplWh4NMNGm1PU7jQUsoVTBal/NL/NM7gr8Umg1j5R+3ERxQzrEcTQl0LLPjw1KNqjwl5kuB1rui
dYyG7Gb1MY/dTR/UIJoxxRp+tBYZ042f3w3CIxFy6Ah84YIKIS4laowwh+SYx+bSqF5mXq1dcp/v
//24m9TmIN5dmvZBN3xPE83PE1QLZEhVfj4AFaZS/N196jHhKfwRHXJfg/JPj6AvOtDRS4dtr69P
IF5T3VsHOGl/scqngLpRP7RVTbO3TQNzL6Si0HvokNh7q2gCxPXO3l1soN1QmlquTPeuaXiAw0d5
jH82OPr5xvE5oba+NvuBBN/faglpnFaScjjJ59fL6+XS10pDsC1Zogx9zJc2cyFhUZwfdj3l1smY
OYg+lMGjZd2F3HbDpwGrHTMzxHBJ3fGlZMj2cFQxobx0REGGgBAet7gfHyix+GJTzCF65eQt5Tja
SZUk+mr0ULZUwqQbz6ymHhBKT+Tv5sMpCkuHwSPJ0SlwqyblvtnHNQCgoT8t2GfzKPotTzDjE13C
zzr7asL8oDGWimEGFjvvJbsqSrfN5+Zmx7PXUJFhxF1ApfjiWtbvbPIhJctyPlYqUPzrRzThgo2z
VVW+djlkrOnRj/pJqoRI7Swn7Vau3ZmVSyvRUgtpCGBSTBwq7GYyWrk/+DdTaFgKOZLOn/eFaejd
IYmzur8C0cYEAR2ft1bWM69nrGxLgDmXNm0GXW/FaDwaPyi6jTvnBlWWChh1xpm2sNCiOmUxOB5Z
xcHLvu2zzl/YL3x3VklQx/S0SRNRYgRv48RVpHK6HtQd/pHY3+Pyl47draYBvnfrOjUxHxqgYFgE
fnxHGblHh1lFG+t/APGKA1kJ7ZwjOD2Pe6AgrgDKJhlxrGfZ5F/MfYV1yjYsE9D+koW8lrBT5lDh
y0hMOV7zdGMYQaZe5OK4wnELtuo4qlVnihK/oWo8hauA2TTd14mZ9TXoOtbA4hoNYptYzuvx02th
EBROtsqGzaZgMvuS22orEBgcErIiCLc7Qt+rr2xiOhOUniXldbANgR+6BElmjwhWyHl/qRI/R4Zb
3CUsS+abjq+yXlKSTpVfyAOHNolSNKU9xDusGyTLV+wA3RzYg6bjW9FWQ2xJHoHkjesLz/ej1J2x
Gh/7tfyeJFOUa/hMrPiuE+gOVyL/P8YjT5bj1Fy0GH1P3qsKlW235CZ/bIHTzmxDTREieNyUyE+x
dPNdBGMvC3as5o3jjDwGALFBhITTlbuIAyIEZ2Sr7v5EvGjBmGWapCXByE9i+6B/m+EmWm4fo/VO
hYdwxFjfWBDevqYecbg2koA8a+UIv9FIJFjCbN4xehUsEZFyapVF89fqWAC0V+e5fw+lNk0fve92
V+fefcCV45kFVM45nERhSBYn8IakZ72xUqNhBQsIW/mUdFD/mNhLKHUx4P9QosCGIbAoO5T3+D8C
dUgUxmG8DYi4Mum+xwqyD19uteyVrI2gPyvVCvhWq6P5GJzpSdN9Ih6bjJgrmpCBLAxv3PqOOMpZ
Uc/mBrQlno7mWpcuK+QBa8/W8fs2s1f1GSxhy3KLdgH6SmHNVD4iR5M9CwHTFYELvQa6cke6c3uN
Yr0t6TAVFhj60ahZjFMJIDfjasIhqGd/aCUcFElQke5F2zV6ZCiiyzWWtVBxQHGDJUMv9pnffBwd
vCgcDYQknmrnx7dSqzGlC5SsLSJ39++WjIED8/hjfIFIKBHjPOEQnuchWxoWtYL8xjHlM4dRWHU0
a1Ga77wEeF2BWdn2qQhIYjGz+73IeINPuaFwMw5uKyx2lWJWHBVTknKAIL/mrEY8Z4jMwlVhOlDP
83/G2A8Fvnnpr1BGkP/QhbRNjofEUhcYrAvsIaWLKGeueAhRFA1M0/fKtbGJJbySya1+xGNN7wV6
S+FFFk+ifocOuAg6qRVZLi8mY8hM18NGc3ZzkkBCmsMADd7b0aXqu78rwziaOwH3cnPoB3fRzOqw
CQCVctQmBUZQersu1NdAqMfhDdtJPgRmFdIFsm/prPg/0Rjeu/SCKdBJjbkLpffQuDRszz21p9vB
IC61mtP3PcejW8KU/b16QM8Za9IJrYIRBJJZuM/KAMZsJkSsmNszjpjvwSlNT+CPWhfZIIzCU7wq
pE/R6Me6JfcJEK/AaY2aKzZy5MX1Eo0WbbE1FW6x77iRhzSebutahJjhmk+p3RhS1A6GbultISBT
3hfslTX0U7SWNvWym/gNRQ8w+0xxKYGsnrdzcnx+28Q2W4hJ0jZLzkKD/66aB0mHgL6HZnwKb/0v
TqiWLrCK+jGrmR/xqIQtwrXgdf0Hd1jYQzy6b1IdbA+adi4SX4gXsD7YkPPsGHvcu/QHlxdPHQc6
3K+x6pvFfjrPsjuTNsOX3JpQl49hhXaWIOmjKc1FXMXmaSPUzev8hcetF3umULS1ZzH6SVT6HnRr
D7+NZ6hlHls1oLZOGz3cDHwuFfPkMpuLvLtakZQcCn8IU5i0c4to+8R4HZA3TbUudG3OPRHNE76F
ApUCM329efn20bpb1FYgrCIEo2RqLns85r1/ca76GRsmd5J7yULB9ZSWLGO/O9ZuCVIGZhsFblCt
7jAERGMUgvtUn4lErSpafw/AcBWupy9wUXC83DIJoRqkKv9Ysdkdof75l5fJpfTODu/PwJ4VOR3W
fOf9VrR5LHEgxhvrECeU9VSipItWZAhFiCwKXJKJhP5+rLb2mXbE1CQfgktGTM3VaAnGPaSvZTnz
UclRb72a5CYoQHLbIHgpaSmBqkDBmp/wfQqsLRqZcNEAwQ/QNMussSmT7YS6bjSsKfv1b5cmXWnw
5nJQQpm3IwzSVOAlgHE//1kwmTDUhx5yvPAhLIO1ZGQ0hpUnwcEmy8qwyrReUsJxsD9anUoQhHpj
OPUncZsroZxxjvOxHqALYFvjgou5gOl6rSPT5wEoIuRyXoNNeU7r9b8XHijTpeikxJHFvQDcqyvu
WEasiCUWUHoYh+R/nWsA0JRp9r41XLBK7Ope+pFDvnq6gcWhSv8CP7wdg7akBn+XSW4lUnLh/NjX
EusxE6wLRoQw7Bh3mmw1Vgm2MPXB9V0ai/prWe0ofc68ZIfKppW2/fMSZrBVRPekyerzgjYIZ4pB
dd8h6t9Mq0kMwAXX7mwyAA0II86klT00QK9lbEp2okPjb6KHa0fmS3ZlX6fm6v3cpG2OfGonqhbE
eVZhSuMSsiRNnfrRqxmmxO/e+J8pHKvUHGpWkEL+pJiNBGeSl7HpI3W2hW3+fBTfgJKXlSt+z4lV
DMof40dpCdD+or9un/a1MzOrStcPekqeb7I9zdLcxta/aDHfCDBQXo323YKKUaIjiQiVyfLIMpuD
SW8MxoMontEUMoeYwKs0PgkKvOER5QCnKgnB8JUAjzyg82wsOWVicFGYBirEaFE5AStKbtQ1OVMs
5opxUTG1yItZN+sQu/plUlvAhA6Fy1476Pm6mb6SVYscD6jxggY1LGpIsWgYhm2FJ7qvHS20iyVP
y9XMLK1Oji8/DahoIPidxurkYfWfUgq2HJSwflVC8PTT15PtpXCvxYnE9376r0VUSnmmUpGCnwsZ
i/nmpDCwpzNDjo+CNDOLEIqboKhk/z3blC6qmFFkpzNpGUPkox0DCn3LPKGBNES2gkvkeRA4NS12
chPAgzq5vqxb5l1Y1kP1RLgvdamMbBw2IYFPVs1YoTEHp6H4CJQfpOh6YD0DRYYyx/XzDnzuFgZH
tEHLDlP7hYjzav/7ltmRk+8RsRvAn8FqXwJB4N6rnesA7pSDz2oAzP4Eoge/8AEz9S6Nnnmd4X6e
zETmThug2XKk4glj4Oyd5bfbem+9l0v35O+6IZNlUISJK3s0H6ho4oIsL7uhj+pKyKdOyNIkjoQt
TI6hObIwwLBXywTb2V8GZAIrMJt3Vj0LLwNVmKbbeB3HqLp+EbRCMcQikWpSbR4ATJj2tqB9LU17
Xhd9WkxQ560dk7muO1BkbJnfYKruoXCw3EUebcSAKBYqziMSYiq0H4ZUW+BFnlOxU21VBNaifQDL
q4eW13b8X8u7A52MyUmS6dKuq9VPYiLanKF4xJ4wT2/IpeYkFUwJPic8CBJI3HR/upqE4+Z69AyL
av1sSGsmJQcHXeagycbq/wf77HjCEslN61ArR30He0xsL6o4XiXAHPIULdsbFZdSw4p+8LQvquGm
fThkgftkrXCQyBvzZ/ruUgQ1s5RGZYWkhfmbt19MIqknsuGpaBI+0a0BSe+n7vZfj6n5pHN83ae4
T10GfLuhSIqphweDuwoTuoDPWZG39VbXyxNhBIpoOwhRVq8QyX8+5QDPkCVLPOPgsMV1PNDicygk
jf2WkMivKgtmOxK6tqJKf7LV8CaKV+sa4AYjlYXf/1P8d/2jIbc+ccaJvkz2FluhuKZFV28vYeFL
WzTtEBa9snynwzNb73NPeK1GYsLbaRUqh/fx9zpM/QoAzcPCOvXXVTX23SCKcVYSU1QfIEZf2srx
t5QK12w2OronbM7OBJqfDzpvAAiS0/qj1iAgXA2Gg5hrybETZf60RYKUEU8BVcOW6B2EOBp5A1kK
cvCKkm3C507DA0/kMymj+rulh5UWczcVJNinLlJD9Fg/FUZj0F5/ARAUx5q0vZuH8QygzQCrPFBn
ts2Z51AQ3Usty5whUPFSXMoH0GoAR6QQuxn4vjXEKaaoi2nGrpn+EyZFmj/AYKmjOWdKxn7rcj/t
T5mXsFtlccIrCaVgDeaOQw0/cZz+qFzTmDn8lr2lqoWLEUtJ/8JepAmG2pnsUB2rP5zQZ724jg7J
Jeh75rmSPQ2sXbQ+af2swa1EnDfwfiwlLDvoabNW+X3yAjY/MwaF4xeAK/nShtfwKEaL+GD7DuXf
1zh5yZ9AOTC/1kLPNYBervLcZjPoAftSnk2NNGZLo4hAemljKRO2t5fczSsteHAS0ayKPYfuszCi
Accg+0QeA8UALc0XVoGmZcC4/XJzZ/AR3NCtxZNCW7XcrULOa5YjCqdIZTl14IiRmGtx+FPQ1cfy
iOIRTh4rnybv78F0gT0i+gaSfO1h5FkGkaRbRlxcjsNAWJSKNUDKYXHzTkZrFnkHj58a5RdSf42V
zHMuVN6WuykfNc3gYBJJYYo/Wn/T5q2wS7yrcHVXNIbLpCZh7VSBCyWAGuwgegTAObODTVzDN25W
ocrRWSc//qUnzTy1+gtnbeaBnWSkkpsJtZMJi2lk95Zuc1TeO0Uo6OB4uQkRkN7Kdcl39Qa39fBQ
VX27pUXz3dzUiG3xo9yhnp5oEr4H4XVc8o6MazWrZUtRxUjGKamD1QKadYNi8kvsj2ered85MZie
VkRRhdpqTFgI8dxXogqrIWZohkmKRiK/18qhOxBqJdmo0gUbUYfzAwRK0U7t4QGgt6QaaL3zNhoL
b+D4WofGoCBjt8CPuIup4u3kuD37p+dKwsT//caxzolrFYG/XJZ6MZmYOH/OxLtFzYXRnSW3VLTE
H9OG7CT7a78vZgod+00FzAvOHXfqbUAEjcaGAWnaXoAqZiqYog5vchBTW53CnUU8TTQCWpdN5G3S
me9LH9pOJa+90FBbBLv3kQLe+tumCoeBGxL773Vm15gM/f5CwZJ5+m7ZZ6u+0tknIYDrcAjr+hNe
d7IWxyYW/m+TlnTfYlRHwXa31tXRwSuO4qaKNSilu0JmpJxeBJzEe+aoNk6qtaU4kr7pm3gQPlnw
AbbH9shrpJkxB2TkNMkgcRWF91Zzc3BweqYJiIeVG6hmwEtvkaP8V6gRE8vVNqqYxdQTuPrPBnp9
WoFJBe4W7JoagPAGfEHP7uXffxt7i6WccSZUV1MXFnIjLT82j3DiobOE15NbBqEYPIKNvqCj71A0
Fj25drOfZYgoYGmJH1mYBYs+SwXWbD0pIkfgYKufKwgfdTOWA04S60TmxFkt6uAT9nNhXXDk4s80
pBj/CFcdp/kYBBOZTM3jaAENWFF15TOqxVNRfZvvCcD3nq+up9bfZc+y0SRDGTj4H+asNaVrUjPY
CPz5NWuU7TeyfXCwS4DEOHZG2B9/8Et2mvDAPOcYCOkCZPJZjKnhc8poJW+0o4zYhNb9PvCOED3d
pLmDDzd/YcUrhzOZwEjayfscUP5UDKZh6CBahEuIvEr2ouPdtG+ROaPus8c6owNZt0ZaYiNdU1sW
F286KdOjAnvwdCmPLsYXmVy7NjwcYfvSJAEno/H0BCT81Q9QuIob6m/7cF43cY/2nVYCD9udA46c
FXfCIBY/yAwW5MuXr/vRkxlmipoph/i5c2DnJvBcYF6SFxCh8WvaJ9pHBxz9GAGXDZIKwVjgrxBY
0EQqfbSVQqjJRoeqhbjLAFX30u1w262LBRLDiF8H/MFbtvGAdm3G7Ox0FMwCua2Kyq+LA+CsWa4p
SE9Ccgd7tVjAMDLiasGfiifo84odifype540itd1yokfSjT71JZ8JHc2oIwG+HPbl9tMrLypl2GP
U6e/A6jz+Mc88da8LTo490eBmsNgoJvCZTgD1S6qv9g+C+OVM/ewobwxhFHp5ETzUYuWtEEvN11F
CMVAg0O058BHZiXxHIws0MCuwYNpXvI8fmLEc4Chp0xTD5nELK073ZrZRE/A4ob+lfGrGzhmTV3z
IDESFlBKT5deYHv5L/zahOCxgTNo/1ENlDNtdb7366jr2fDZNjCYaB6cKLqyHa4yuTlWU/preqo0
Ua1emseYUgRJIn2O4mC/aq3jgiP2EYmBBeZNJuYtDvyTa+K22s21U1gPN0l44YvKfO3a+dBeuhT7
p0BWQQ6bpu3SJMeToH63+ADQSOjvTfeEkOSXUJNXoHE9wsNwDzb+l2r/CF1U0g5or2HDh+F32drv
LlGFiQRZx8+N6RNZtpKvCYYBum3uvqGhqGYuB/sRF3BfqSdMwPveRR6Ry3gNO/gI+FPokYwET9WD
aeNEVtDYEmGVN7fR2xiRc349TEwEAxNfKr8Juwi6oPjaceJO/zKTiD6zAZkEXySnwHcPfdiseRep
qB/hSgTq0Jx34208QczTKRudd+AUXuYfVXHUfjztcok60/BEu0xwMcNExjr5QgWybdKlBPKGtLJ1
vKjCTdni/Wh8adJRC2JJtj42doT2C2sGEy36eOtq9Y09ZwqdYORWmh5YWugbKdde1lfnY2WnVSfG
4Aq2awKScOUVzYsYT2ZsrU9XzGsBNUQT3LtP/tAkFxVCTIHgj/wtrkoK1MAqEMe9Ucm7FneSvQdE
60yBejnLc3NxKrsLvjNJQniS7YBLKiAXKOfbuxHRLUngMI6QZLCpaCW9+X/cNBXe3hDUXSMnF2v8
pAXPuOvLl/DS4JXtOD2qO3CvZlwEpPEOQGVrBMFFhWu4uaKvHj3mJPatMqnl07b90um2i5BynPC0
l75VaosTXAmUESIGHVqXD+Xw21jVrpkQdKvtA2y5VbncINpZ0Mkp99VLvNEhTMUqdzBQIP6hg84j
gy/E+8qTvM9eIP6cyQ7VfZ/PtWZcJKRcbJ78/wyDmmNU9Imo0K1fMYCmWlmRnjNWKGQ7c5U4sUdG
bR4YVAm6enXP640/jKMb6ZSr9Z8XIpgmVItnfWP0wzC6HfHnAwcnhfuQ6O+AFrC/JPLoKOwBid2g
cpYd9e4FZjlvjMp8yI85Egzg6xdYBh9HHZksH1Eq1dfcNnxvindvEWljQZBvydYYqx3K/xsLK8hb
49daw3rUiXpTy93wtaoJ0fJx5JhRDBPbN7aXUKdgzUBZJuV2EG4E0RKoxKclBP+TJmsi/T9CP0Nf
C2cYqtsegg2spZvki1MBARtSHctM8XLrp/bekGW6EevegBDeFNyXp71lEgU2OMvuG3R4DMobjCFi
+oEfYVs+2FgfmWnPHFgw4/+CaeF1jw8jp1Qi5tXASmXqCoj6tHHTq6Msf+aQN+GCjIaN3WJsHdu9
RLNtd2cAustU0wAC+gJ6USk1p+jvKEBKYOME1kd13CMco2wqHzg8v50OeD30sAEYuNZqVxniC0ON
OOcN+6Lvwk0V0WixnMEOo7j1ND7zF1lyuYEu5CKYqahUfO0p0uHGrNmqMoLoplQ+SiumRqqsuEyN
weFvStJ4ezCLYjX8DV7Ok211QyuPhL51+6KhTEAXHlb24pLWlQ7CITl6pRJPCf8OXDSRsCHUbKjr
NBJruLUSJb2COcxumXs1ISdDnRf/jlLNKKFbAhqS089Hr+EMygEQaGQdF8aEo1UWJ0a/xV1UkULq
o69o9oVSwdA2iti5qncH2gORnSX7xmZmpU28jdvLcrT/yGgajFpQOrKvgh74lUZE087T1bJo2S6q
SXceNd2vZiZYYsIxvD5lawVqtcGHrD7qeXr+MS7FwTvLrL+zW5EvjiWnocs1Jwb8ph1llEdd5S6G
oMgMFFWvqGsH0PhSUU1ghRQ8yaAIUIqkP1SA6WYFnlI2I0NZiQXrZZ5klidxzxXSw+SDHaGIJqwW
Xy+ETEjsgSMluYt4Qhf1VSQzYaEJoFPEbmB+i8TtbZKYEYKdjskVQoBYl85NwS4eb29P6Bi4kOe5
E7+mv7pKFldX/MDkv5kzklUZJANXK13pCkSlEK+DHcJDaI35lUg13jkKpL8tPlDxcQBYkH32VwpK
A7iuh7toxH7V9mXOJ7sfKu+u/A1PLYsOjMnLQQb8mlgINO6D0wUmVbvDeWAZ5cYi/1o5MJa3+uJR
BNzJ7+g/Jr8q/I63bfcvnUfS1lVX+52H5OEfl4WDTLfe4m76vfM4dmyr98pum2E+XW5W/5isuiR0
uQLSwI8zU6D0gBOqoImVSVlZhDbqXKUQ3GTeRxkW44iYTIWbdYigFMXxehuO3ef4PMrlWOnFofqg
+NLMR8E5lU2t7T1lt6NZddcg1Fe5dXsAEBN4onHWhi1XyprlFQdjsu3WynwZHF6CBSlb7CMLYSaQ
SslLdgfoqIYUKG4K1kBOmillCWO9gKA1z3zu9Jw0wsLjh01+cqbtrNIYSyypsyrgGwWNSDsNVVA6
1iXsfYG06uhO22xG+stNEMtGBb5W0+Srm1ZMHal2aIkoIRfKOTxiuVFCWrGZPkuH+Jd/aF1etdwq
HODcMKA26CqUESFbwJq+c9OIGfbnM2NwFVnhHuIuvRUspX+KK+DLxDGqKp5SQlW9xOBf4KVuctPg
62sU0YXFwDSvR8CXXhD5x8BBC8RggLUXw776oCxULnh5+xOCMdVy9VQWhVugpt3t85O4YPeGlVPM
mxuuIRI4Ek9vwntYr3kl5VatJnexVLJ2oT0Q+OAtkI8pAbk1dgoX+w5pWYl5/3YCuWbE6QjqiL6G
ue8jNNXJacdyTiHx1TraK1KI4itFuO6ANDVFr3P8TBCt5ds+5a4JsbGRUzmuK8RSQtWrKxZ0Pk73
3fV5vJo/Y1iR6c1ZonzoKaf4jjzpilbOCYKzQ/jRgReAkZcqIOp87FQpfoYWYNVNrmfQAvnXqUZp
oqRxyCsdKz6Jkw5Bx/VLvnFrIKI1obEXSRn0CPkWYDDqwVdFp1M8IzYl6UB2pg2G7yURjJ38KXFs
LaOwY+jyjK7aOjlLToN899fu6rx4Nd7/3NXB/aoDReyeB8WBcm5CosXXxAzkQ8ZJoCa2z/cspMLL
KwyTfWuNhcA4O8sTafHyU1RKtx+LuLmVYvxWWRrhXl/FwlRG4N0sp+R0HueW8BGvCMg6n8cBg9Ec
z7fe0DrhwYAnFQ6MYEBPyWHIHGsG2LlA1y95FONqNsGkEEPyAUW9FP28H1/R2+lNY+40Na7erfVx
WwqqDL1PQHOaB/nOk5/LiOQ0aXKtqUlA8HsVsqp3XcB3LnLAlFa4stVO2viFNHCtbu4JwMELlSvc
c78LYtclj7l+8UhlOPwcWIbnTABGdlkAGSzWRQxYC3+wxZcvjlVi5ru1ampFWzHlwagF+Q5W75ap
jrWt5pK/k3UmFPQUX5l0G6WWhqPcf38mV+pOvx1rDN4aCocucupvyn3j9G0JWJav2NWEaBqJlUKS
aqmXIdLpFDRtkkNiqaBLkIarFgQiHHhy/cs9CvVkvcP12S+N3BEVAqYU5kH+2HgBPL7kr5d4sPvR
r6K7VIRdjNlnSyv5jhF+nhwunul52Rp/qhE7ZeSs0HVPPCCaDIIS5/Cke8RPlc7p3EI+2O7o5c5O
8NBEDCjjokisXJX4N2h91RHFwUl4MQcd7IEoyyM2X6G1ymQuhwQ5uPMC4FLnKGz3FqWrzPKU2nXG
XwlFaifKqD+OvX1fFbEnNJdux7quX51TMiOBfFa4hYzcV0TKVL4KIvcEvAf6DS1aSvCy4WBFbydm
13MjvQVfydX81aAl/MnH7ImXgV/sofKhK1I3KK6YMUu83Uu9X+KearSOIAM27ZwMowcJWCpR2O3E
KpGLstEltor7EKwP+QijM9NEN38nXz1WF6nJpH9quuLWA1dYUjz0ndsgXSwOSpK3ZjEGja37sTMS
mCh0fS6Q96uH/AwHpeSIC5ACDtfZzbZMZui9i5TkFVU4TcXSXGu+wAarZqwZ5PB5yt+wc+VBatIP
NsrlaOcPS8xbDq62Ajrg7Bse1PtI0ZlmVQad6gkcW3l84cu0K1g+pie1VKRzVAEsegjea0JKAoUB
Okkpb+xKKQzFpfk5xL6aw+jfnn4b8OKTYBFIR1xoEZCQoXEUhNCX4+KQo20uvJ+weEjw/h9cvA7w
K8vHuy5KPW4MLhSzq0F5w1a64gu1rsWWpTaUFkgJa8jjlf8laQYHvvDcjvUJC88kP1Y3tr+an8Wz
VeWDI7NoH43wuhPhuX7QCPQek0VGUQdFeTeVvSfRAJrwhHLmHbWgnx2SaGwdLXjSNwodLgbjdAS9
AgeLtslO60oiPPSJMg93RGU6ubFqrvrFAa3kgaRS03n4iKuGxNOh+3h8vvmOuH/U23tFCIN8Lysl
6msFrpf1AG00JZIofgAtj/VvyTOqRbO/tKvt9fUCU5zHI4VkPC/lpOIuGX8oYZp1hdcy8KL6Hh4I
gFMhI8CDA1DbsChBwQW6+XVLYzuJsPrAayyQNQ/R6d7DCgPLmwNqA/57hdTuxK+sJJA8G7kIhlhH
56OmIuvcW5v0+S89jTt4UMqkTSD4Bc8BcfGe6A9pxSApRllyXIbg3/hjtYNI7Cd0ZkzAlt1R0xBu
6ediUJrmNxHRFEjDQOex+7rkvK0DlBxtIrtd54D/K2P4lsIV10yXZOuHoQrRMrQ26y0E5E9IX9hJ
FBAKUfK1ltcvxbPUOtrjPCtoRbRA0dF35itXeQQ6x+GVyc1NtTwWBg1ylh9cLxYemMDA8WZ1CNgq
/USXXvo3k84zpY+fPUEMcmGF3bJG3tQQBtRWD+XofBogaLv8b9gIPkba8Ts2LjHu4Be9Eu7BZyLy
uKEoLH4T4x3rRCq/I+bdoyY5imEGQZKsdP7bhGA7LN1HZEmjVKQY3HYuf8o0arXQ1nwuNBDPaSLY
jVfl6zHlWVl3mJ3YWrLvWiQQ1xeBVcHswATaKTQ7yfg3DRk52bKBaMOKUqCqeem9yESxvUHioTtM
1uqaIrwKjojah6kiwOsqz/caMFWFmLWgHNPW+Ct763qEBbY2NnEx3bUW12qVJ/YEAcWkiYg9jbfy
GDyns3DT0IBxrwleiMQNfqSS94phQItFCttEDJQ+M0fAAtaMABpheej2uRalTY5Mj767/9VQxzHG
QTrVU9ZolPfdEq6lc/t/3fSSDAdduwGu2WqKyR4oEkwPbcDwpFbIXI6Ndehx1VKDurSbA2GGqr5Q
nWRTZI74gfxoD1z4VEqvq5mC2+eMOTKMFFF3cRucQV3x1jTaVLGG48l+pnCnBZ25pnp3r0URLQ/B
SdaQbbgBGYMHJbdCVuMCtTkvXz4Yu5ead92oTQr4g0fiB3ovEbxlAbwijIBoqAqG8GAcrH5a5SCV
II0FUKrGb2lvTjrSff6Uq/kQixIKXTjjjaeTbwAKu2mao8YLDVTolzyBvniUe0zkqCUB0HJgYLfu
H0+uwOgFHITXo3opvDNuzAM2j8a7cOhFkZm/R4gmIJyPFG+Hi6MVxLYqz2Ah/rVl4YAYVPCso0Gd
QwaX04EaP97rBHNJNU2UUugtJ95sn2uasPOEDAqJNO6au4+S7iqcvzP+7CA+42DSK+8RuDgEwlas
kUa07Ds2HUJwUJWaoHYVY1uBmdQKdNWJD9xedao58R96J3Zj1D5TIsMjlSwTgRNJ2J3C+jAcHr4S
otv906qZKvNTqJYrvOzJHpFIcmsjkO+TUXSJuj5M3NrH52ZXGiglcJvGjfc2y/1W2/6LwGb3PkIE
Uj3g6jv9PiPPjmCk7xsgTUCYxQcTLbOQ7rbfwIKZHGukus7vYKCLM3DxiaMpjrby4umOT2F6+FBt
mieeOroVa6FUIipWRVqoiGVLtOKCdj7BEplHDdeMpUO+eQR/oQFiC0qCA0OTj6qpXEtKsunsQnK3
CU7cpPD+GaCg9zd+XCEDQ7TRFMDXyerC7Bc6yrKEM9XHKRKQDOzMFpIkFpPWbdHXZSrnPZELlQIS
YOTLfLb9JkvYPj45S7cRe3qJBX1Lg/tU+O0QJnAFGin4zlJKtD2Lp/GuIOsgnnkUHyMvSuqa0reg
r1MuTSdkOcKKHqqbD50uxoRVWLlmiaZLYD9rQtSiUZFxW+OiyV6FWmIzD5qFb19iawF7ztThapsB
0iioQDgWLplcwrvFbLHD0n44oHqiRkXjoOxDzU8t6t0OBrZ4q0x+kIpPjGoXB33yRphLqI667vIj
aHOTt7UJO4dqPchUQgnT0tadJ2n+Yp6GWeEFr/aKRVWZNWaf5i2uyX8EGINJSxR++JC2NBxx6+uP
SVsClPj0OzfXGIHmMpEPu2RMqjUfJtW0vLrTs8/0aTYgo5M0nzRuU/LjzYY5b5comJc68OrUd8r3
cDHeiwW9cLcUIZMW0MmkSxQ2MJgk8Vk9qkzjPIYeJGoOmo7ne6zEr7/lErF7cOcU1PcnhCx81nBL
evVlWIt6146o7ZTWw/TChHmgjOCpgwNj2iEMA74S1gtu4MHKKZUd2tGHyU9+0s6clMPPLJ4znZ0h
EyxKGtM/EnpK1Wtyvntz8XwH4C3povX4rQASI96LsBrTXz9Us6hf2l1arDHI1HJ41yJICJX8tl1a
ZZHJQF/EFLoQnzAF8Fl7R5YF5iIvGCoMO49mP4WckA/V6B3e5Rs0hzmMgFfqqmv9Z72KOyOLGG8G
lb1IAgkL3QDWRl7/UdlIuZ1HJKDn+07Iepa2B8Ef4iJo+PffsVbRnFPa/fjVAnMU4l5Ex2iOvhGS
YxnAuJZVCp0xoBjcsatvaMoF5aZqNE7fsnyoBDQyyr9ZoEfg9eN2otuuz4Abccug3AV/m4vA+7j+
2zk7TW4mXbaoU4baurnLUtEOBFCCYyycJIwvwAY1Vx1xaj4OlakxE3x4z0mawaxtJnrS4+jKLS+0
6P8bs4+zcUzRErPoscgvdepdDg7czsPQU8BMbgg3S4fk6FpUW1/KcU+oTVPYxjRJ33lk2HzoAjZg
YuPOT+syklqCAtLR4vD38Vmi8jWD6F1Pifg59n31xUBZQX4Be06UieYOCj+Nntt+BH1TrhHObBMp
7b2aE+AJWGvL67ieZ1GOay+ryGzYM7BByTLwS3IXQC7OWyY+xKh+kG5j9Gp9s50YzrCKNOX0p0SC
yx4FPhXhTAiIztGceOqXs8DB9nd8MChJ8wn9qigavaXDkd4W/Cm1pmbSEkRVnpZb2p48uIe0pIlw
limCwzRYDvgf1h6lLlMZDWEzr1JT07YxPyLGtiwxXRo3d1lOkfOZ8B7EVj3uHY33M7cpMdvE5yJf
IAOwdegP3AQAbucxTPx+/P3zQj93XUNZngmAHM/dmWffYMuJVmCMcRxvSva/g2+lxO9XeX5qVIvL
7nWn0fO9js/nBlMnwUDvsihDgkgUik5ARzUKpes8w1igLFx4ClmZEnGrci6NLTGRyj2s1XB2YcV7
DXu79QpZDCFP9YQoQoBTmN9pyCs+hD9msS1Mb+moNPmucDGlImA6njHUNtYAyQ7OI/QKymqog26/
XNibSBv82VpUtKTqgq5GvbWAHrp7S1cchnzcai1GsoLEpa8lez1eUfWeyZoCe8rBQ+7BOR4Wa0HV
sdvOx9R7Vs3sAH6F/2qm0RKQ2CaZiUIaXj+hgPWGIwhimJSXSj7+bZpD/3H50RAwTsUug0OYtf4G
eEvFWq0mDp017dZJRPtMPoC1rzhn0FuR/3MOo10JTAk77GokouRz0XGIbBtzDWCW0PE2r32U+PSU
NhK6fbBwDIQ/BXCulhC+fU47sd0Vd5OLjVfNj6NCseegQkQhfHSyvqoYXTeF2HQUflEfaerZH2az
EZqwafaxV3owWGsEuLYf83kTT3cePtJXBzVvw1ZMbX4F1Czx6SYSisbAlH35HbWcmgZ7xhf7PEGW
mv9LqLsUz/U/93ZfPkILV55+g3a3N1XuhgbpOtTRvhWMYnihNI3eNyw+DkthMHVagDI707ksNUvR
swqOk3Lv+BobF0WpAu6imXU1oe12vULFpU51ynNHMeGk+ypbB9U8utoWGOh1ZIdcJn4Zs7le/G3s
uPDLs44imXqi8421pBYnDgx/Uro1IOgLr+RooXGeGlP2uq+RRvNftWS4W5vKSQ1E8unw0pPH3d/n
yiPOVh5R2yaBDZD/nIP0EZLhwmSQ36ing91CGaIJjD6zlQK3KECbtUbqOcJ3YVZ9c9utvmCjg2zz
x9qzRHr3knSWELhjD4EFxoQQHmwJPtbpan3JqjElU7z/f8o/JxyJ7ZFY4/PqR9d4NxcQkkAV2GzZ
0gGO7q7y5H4LY3Bm5krZaWS+sug2jCYvzgxxRaxy9ZAkOUmvdvPiMGlTVAQv9mxweJYrzZISR+0i
MlAXvbRjkVDEWs+73o8Lzu6TFWbo+ocbUkex8ESWWUw5Ahc19nFY6I63re9gfbyUe9E61P2Zc++o
n87jvbfDFp72tlcgV4LAnaWysvrdfAQ6IXX2l0Tg/3GxDqxf4/k7QVPKFbIf0dGRGWGHew1D821K
9wmnXNSGLSQnlgc5RdfvBUaxpwJI4T17LcfkHd/xU662kuIKiyA6Cf3SKOeXjcEnF8MnfI4wk6Oa
2EF0azxgN9xL8NuDXVDyLIhb1ljbhM+X4GZaV/AouRBGkXXITa/heEwqX7zWv74ITgFVIrs9F4zB
e3gsGpIQdTY/A7bzF1v3uROjJVIdOdSV/ffsaLekc1obYDyrPq3eroFpujkC5U4JVts6zHau8dhA
YAk5VLkzgLf2A0iHgyEGAf9COd59+so+QRQwPKgdzJoQ8YcKgeU8bLfifpDKMW2BUkmqwSkbWBMz
dTc08mfKZll5la6gI7/6360Ir78Ke9A4axCyRCFL/UjEm/D1fm/bOInIJcsTXmhPI8D66M5bvbIT
BfDzC7BPgN83r3tAwQxD39SidmpFHr9HgLvQr1vW2HJv6uHzVokoWanE7ynON5dkZw3Cz7m8FUXL
6z+UZcrCYjjgPwwCNkzqFi01TEQzAcoeDjcQgKsVZ7MXq8YphYIDXHyI41wK1ug0B6U6WHMMIOMX
4mbfxmrubtF62hB5g56UECk4UjzFqc9lQH9XzWm6+pLzsPLb5byDpKqHlsj4j/KXkisyBi9Daa7P
7tdqDBsy7JPKtcJinVr2IVEgu+lbZWgMzAhxM72oGhV5ynQQnK0Tbzrz1469nkZFS+U1OjHAwn1Q
tVbaECk8Mu6JpaO3kylYMVf+7KbX5T6cpgrbgoWyUWFoSDO1YGX0FKt1CTvlV4xinPRn9LufV11s
cUYqJmwNSy8H7fS2Z7yZCFwkepM6egSX1tRrE5S0nm6ef0UkWf3K1sFOUMXXZLuFiAJjJvPEe0Hn
jx7Wr7/is3Yu/CjxaJHIu7DiaSbo9BrFuapdcn4hbBhRJysuUh6V+2o9gCWsA53oUDLlYSq/J1sJ
3Q3skvvzGRQfazlHbCYwJ3zcO/7M52ZlUnoyfe02UBCnaZrYfQPz9qgCQyfCPNY+qQriw3BAT25S
oIMKRP5EKQEsXldjp3PodYCREBZGV9sQgK5wjFGnT35LrCSfcw72aNg8/efPei/8z+u32wLJXrpT
6hZVX3yKNBvBu8jwat8wWWBMsv3430fOV+7xU8JYe2OtjBwTi5rlp3zS+KflYViJrTYAyACCnMMM
la9cHpH1G6mM0Zn5dtkv2DUEwqSOGIKc7SxKy1qMqBMCNXgYOPDr2kDmSSFuCekE+fwCSEUV5UT2
foIbRaTB0pRR9CI073BUHFv8O13+rL6yY+BhlT5g7QLX3nO13gddt0Q+AsaqO1Mz8FQ3cIaC8rzV
mq4wNLLrY6z+Z5JrrJ0qlWUh7FhPdK9XyHQCukBKIbulCHDUe7jMNOqSFdb1RvEimfhVIuZ1c3/u
P4GeuwY98mMBrl37qPkDY3CV0BHq2zweZiOsPSs5oAuz32zoM7no1x7Hhr+Er+8nYwXHIMdn3Llo
6PjTMeFKJE7HSPIxvQmgWO1Nf8hsuWNnpiGcthEp6LMiAYebAFxIJouL1TIp3dUQVjfOBLTDOMPZ
k0jWYikKceTNrHNxveq+3Ft342BPXgonAmVkXBylqT7obplZi8nfCZ2ZoeF/68VVJ+tYGdmM601Q
DMtD6v57GvSTZQi9Y15So/PH3DBxO3/C64frNdR8U+47KrnsQst8UYNW7+LHYq45qCfnUCeNp9dO
r5rSmYo/J0Aug6FCscwqNAPwh6h8TKn9pZSaqigTSvsNJfjbEygQ4xZDiYjSI9ymFp3uaxx6hRg+
CWbBnaSOEQ5WCvvtEckcx6BgZAwTA3EPi9su0i5yPHIZcTket3f157XuyrhzGbsTkOCeQmEXk+SF
PKDgiBDACs6fvhqWbjBUCnIsROKcVhtgCb2n0osnWczIoDsaXzHoVugAgOugF1WeIP7VC+V2+Nyi
N8Z/5hwa0ntgwYK7dLp0ji0a4aIIXbGu6s9Yk2YCJrFvdOKtdHyuVu4vn8Nx11KOlcxs+/95u+Q5
wzYn/WExgAR7dyJ5qOmZgCscYpVaokbg4Bz6nkaeDeaYc2N8BAceEvAB4L7zB5SMxSBBgaNqk0J6
4Mj65nBYHxge6wHz/XTRWAqpxHPrx4UoYQ1Bjf9CK0a5Yt9lwlCfeTK6o0c9xHVjZlbWMjnckBG1
7SkoE9QJLP9dGZwrmMiOPCDMXudk7MFYdD8v1VOZMt3OsPiEPO0Li1xxp5SWDDTI8kVh7FNS4S/H
3vSwEF+DJbrkq0MZk+5q1l4cqe1xeUKWHddyw2w3tH2L82n1LIYskIFUw9MwUTUN5OaT9dqYMNhK
SI07S0D0Bt5s+H1Rb59lRmkbXBGn5wIgufZGmCdVX9IYn0A4QDassIvU3PYx24CTdvr228EALqzc
3nB9AA+r+/Aa2CVXPYNjik4QHheSZM3LOjdiwLkncJcMf3Un6mEr5jdzyjJeyK4ySn7yVQEydIZv
yvKuPg2gFXb3BGOYM/9jU3WMiMnDq67q4tCnLHVsarcocec/9xAs7gJ1ttvE0pijvJBPE5gsbntW
8v+2HHnos8DAsyCQm/TPMADGk8aC3K9Bv8hweiAFWcrzIyyTqFFSUDXC7d3ssAu1c8yWrmVWPUuj
K6GLd1dpT04pnvI/MUBvAD+OIGdm/xPqD0Or799CiMRk8R1FtaqwejAJJmhFFkPWNBFeMomjzp3w
DcfrJUQCAsMBaINNdWE3UUeGziozomxKjRV09cXm6brDBjBie/BSQvWo5qBWCiTeI7dZYDxC6t55
YLQczCXqt+Y+FQ7CXB+Nk5vAy1iokXEoAhsi3V48kawHX9q2U6TdnvIjoRGwlZ8p615C4UIRYo8A
MtlBaHiCERXuSBJWOaFI5KnhE/i2Z8ePL3l3pHsYtVksPWkS/WJTPkjHpSC0pJ73khD2vZc7B7uQ
w1kbvBvBy0aC3kvOihcgPCJfGiSahIlmcEC/R/ly8A4ZF9e5bebiL6GkYzLkRAqona8SC9cFhvth
Cwx1rmx9ezjpsCQx+kaTgqcxPAhAJAe0r3SACtRjLymVXwR3woXdLh7qJ13xI4V11d3D+xYAtRjC
yoVGdDEjZ38FSXogk1BOt+bVx+6p+LKbz0foYF4Zz1YolRMFdIPWKhDtQxN/NyVe2zprbukvfL/F
Y30gfjFFlJ0m5aGTuK4q2dMBBIyqfobyi9PB2l8Na7dOBo2cL8hb8e/ABs4tCTBR+fc50W5MZy5c
DJ7IhE38O9zTaDDA1u5bK1NIsWmQcY1gbqk80vl23hr9+wbhOqvtE2uYB77Ek/kClPX6YnHPykEx
EnBKpJzYIf2Emsqx5AWKcKGPPI/RGe6jUXnTFppMo242nT5Gz/op82ThDcQqQIqNBNtwbmtrLTVH
AVjFzh8W/9VmtRJEnPmdk7xos9qF4n/FWsxZzytG1FMt/+WdmXNO3OGPdyZtwwlQUyFJEaH8NRR+
9y3M0151NDrk2zZ9uaLiYZzls/ieSeYJQLzAOoONOgxdzHmBlPC8Ph0vsgW5gYOuztnm0n37KflY
6UmUIp2IK/O6Wy08acd4MEHFLw75dv8ZJVuEBhoeEAn71g4Tzu72DbGEcvMwbkSO0nFRVo5bg1vT
4Xd/U22FNuc76yEwf/wybAqJQ1+t/KJT0WW6JIiEB/wRebbgGvNqtxrOb//0DdifM3/DsxogST8F
cFZ5TMWjBiN3tlxG18gYYHfEghUBFAbATjXgGZ0FUp7HeBJgNo49R5jrBtjKGKCX+Llmp7XOFF3e
ZVSDAZJsjzcv/skJSOzju9EXpvhVPjjOUbFXCtx/6XVUCx0EUnaqivWUKGT9BVct5rM2vebaGkxt
GUrXc8F/25HYcYSrlQQCtHUTnH4g1bGwx+qWY9JQKN9MhbCM63YOj7uwbEHy5sDfCo0ygP1Wsy4g
PVUHq1ACffDGvrKed3CI0V75s35oBAjCiO8U8npjWFlc8GcuJs5NPW7lkuKJJYvYvvHFX2mv0hSw
ub4wALe1KWJSCXq7+66ow+dGvYJ0hmtHtyv1R6vc3Yk0E60uggeENwdxtVcVS9X/ifgnSz+0R+Tu
ZdOPzlYbJsEc2jvKrnPNmpMe9sypMBxQX7hCfYGCuaPQnG+X5SNTppuKa2OwZ1afn6tbdYZt/nN5
etU1oDCy4YeLKXTOjoNd0sE3FfoRnW97gFu3RCnRsZNc+Zg35Xb9f8GoZcPW/LxfYdveLO1AEHJj
HFZC4y9JXdToAObcE6aKANK+qNNTs8X4uZBVHK5ZknFPZ786JBiOwXSxx2F8S/RgrOCvpLKw/K24
4QjG/h154tYjImsK4SRq6pBXW26IjPhpJJefCqPLu+wUlcpptrLbKH0CHaFYF8kM0QWyCuCrrNak
ywT2syqPSb6YIVC+0tFOCNLAr0ip6yevgI6XIIFyUo2LyzPtsXW1CjMg8bnBE9bT6Ua/PGSb1X/y
ZKSer9arjz7B3ga3oMg+2crpIcrzmvf+JmRyIYCbNCqYYjHqSANx5o1nZnUdeR5YOybcPfJhXAWe
sKe6gTwPy+dNS1eZlziuDzob7IdVb37SYAedGzctbEgd0mC5/GkjuuUf6gAzYzu1mREKNoqsoSE9
SUBp1/rCAnSGdpXnBKOkOIjbbT35JXKoSOG3nfnH59V3tjK07FESFPBg9CrxA2/aJq8HdnIAYjyb
intzQy7q254Fp4B8XOmT+HJifYvfIPK3Gaz0N91MbkL8I6gL9gjX+r0pHuFYt4YRTvgG1w4T+wQX
PgueXfq8Z/afOJajSfQb8cz8e+iTyxUDL4XwLLGqkzIjKirPdcDzsxOGXE0aCT9eAOSmC/4dLVLy
rAY0n81TJntSy/X0qtto38L9L/0CHJtcT7qmeyJPDAOuJmRcBXw83LpcDoTOIkTy+2P9xN0VpGPG
bXnBeeK8jDGQZSZAEOvp/hFibB+l0l5XInIG6jStsUOWd0Xhk9B0dfNpv1Gn4qBlmjoLfe6ms404
wH47ia95OafJOeKXXAtukBmrfIeOD9R7hXbtoGv3EUFBvB4FU3QAGmQeb+YF9O+JVEuXHvoCVC0I
nYyyNn4Lk+ZIEMflI5qKGAJhi9cchx9KiTqKA6OchQ4xxA6DQf686lLA+m2ZD2K8chj5Z6dvF4KA
C7gz8NOmThWVcHOgWAJ+IK72RutO6Js0mBckP36N/V7lRUwfi++XRPwbRdnCHqCsAcGmvj2ELD2J
0+lbYOv+ES300TISX6/1hMTEtZdjBOVLOa81UAq/UqkrD7XkPR1EsrORxbxanPowTQTICGb+Qsd1
anVB11IFgdBUDOJWrKHi5M9r1UCAV1eoRyYKdf+VYbVsiNLdA7Yy22prN7V3Fy8LRvL2zA/GYRpJ
15v3jzDpxJgz+1fV+OCllRC6fzgT1yZrr96XcopsTfGRNJt6cDO8KBb7UlpZJEpiReYg7TEa0cZY
NuZQIbgNTzW3qgkj2bW/1Tdl+/0kEEliJ3HBKFhtZjg+qavEaTOc0VgL5bL0B5iiHD4aMa5BW18U
Nsn+jxDsVKbz9aORfjcqFGdl4/GaZa7KUV5G3xyTZyMhUowAbgzFQmPEGkumStihOE5FClxU76xA
cD3y82zsHtBPt9hoYC2+FW18PLJ9i1eLI0eNl9lDINq0ozhioHJ6NC3VbD5tLFJZCnLIW2r6XWV8
W0O7jFY9pJ6FtkcCYevZw4XRY8Kz9JpQkuzArAEQLZ1DnBNF+diAqMvSHm0a2JJxeyAJ9feywHgE
06SBHhKbuL6Pg47Ajp8ig8q5IACtkNMEpZe4A4LliuYxDMhy7P51SHLSjVnTKsXfs0wazdpfgKTh
xLWTFNxdN1IHouiFylzT2nj64W2DTAI6N1xypVP4OlAECXguAhuZ+AXw6ZfZDy2uqJOBqiuSozU7
jziJxnYP1erOa52/p5BMCKejK9x+kUjIS/QQ9/qr9wITY6a1B99uy4OBLv4ei/eDCvKogdvQAsCu
QgI2iQbyssNXADhAyqApYjcCXFf65kMui5ztffqCqBK+6GlWAp6VmAzu2sJjyO3B0G8eaN0pig+7
jS8jQdKxyZqDW7jtM4Gmz9rhjtlLipbOLB5OvYCjglfPiN1vkcVEryc9VI0PAiSVIsGuOPIxoJnQ
D57AUlicGQ/YFP0p15XxbMoBAEnJ/DghQ667R+aw1O6lqxB2eiH+Uqe2vcaM6hQN6+fExIyIVFg2
SrzdetECsWLzXNfahK4SlWePqXoxlqswzASO75Z5HfiEMgojhdrZYn6plShAftvzxvO0CfkQzdUa
wuZ/3rVt5VlcKQRr8GR9Tj1CXwTTVUURqq6A1wCPY4g+C3axf2n/Gdb7XRxyCWUFC2t2p0hc0X3o
Cx+PVtQQrGA52eJe1mQ6u5tk7SvJIowveGRyzfzXhMvZKMCs5YF5kSPDPs51KvLqrozv2Nv37m4/
pLFsNjcXcnUPQ8OkBd6h0lYpg30tMmekZLBoJ3eCuXc3DRCqPJ278o/hxPPuc8e9F8NzHtuEJhKR
4zm+6Fiqzh0UnbDnl8WC5ajNfZAsIgWUlH5FdV4WW3DjyplEF0XPOQgexPn/RXeZpczE7IwfSzoz
LtbriqmtglhHRL2Yp4NYU6rYl4ze7fEhzaoft042epPy/FyM8fu05kdJ9UnOUma5ZJOmsetsEjb8
l83sIh1VhDHsLsR3R7/5JcsKvn37/ubA0cIvFa8SDiHzpZS0NSsK/fVAhNzNC7UUiTYAoGnYSJ0W
WIsrBCxIyoTMkZhOfCc6mLRFdZGBHNFC1FFWDdOEoBbfcpce2iOl73YNO4NV6Gnsck/zUnZKrf1h
YtYzm8NA0u40HG1sfV7lCQEWJu5LY4/NNAw9LLRnzxJSt/sDOMTuJehD+SBWeVzsJQ52OZAx+P7o
43Xjm0TXPa4u/Ffa9OILX8dMjmjyPUHQnwrNUxmfbVb3/s2z7sy84kEEAQIQHDEYuqnirYz633xp
/SEnUIv+6PIa+TZpjI18r7unF3uTwbjJlyRVdG1Qp3AY9B+IlB3vusI2fEc09GIggT7Tp6MCMwGn
TX+zym84HPiEkqzVkQx1QsA3BBr6Ja165FQ1reDl/uzXKJEOSjdSkH1ZXvX4kN0LwZa0nrvPrHe8
1xqdMBVY7H5ZkpcVCZVYAFMZitzQK476xLKsvUqJvJj9pTZ54JSxOq87d/f3FpHtdKmlTBwQ6mwp
i5Rj6IfhFpqj2gtdpWsF3D2mEPVKebyJckMU8K5lVUlGk1O4HsHAdkx3rgaP5T0VroIRR9m8Z6Cf
6WRV9DvEWmd6LJg776UGvTJStEFzGwhJFvfFsECWft17+C6INFE86vMO3vjVvRk7tTjlMBCUDCL9
JehdH1/NFsU5AeR+oH+rgsom9k/cb6OI/qDHiIhZ81cKa38UoaQjE8bCvwqpPE/bh5QKsqjbA0Fi
EBxVOhUIsOS856LtU1CjW1HD79N4M5Q03TBUT6dIYZbj6tqErt87fkb0OjUw0HoKSZvrAOzr3FBk
1bkTzdE78kKuHLfFimjuMLh8IUwBPE+Ii4MqmUUksvAyswou1gYpv0z2O8/iPPTXAN0hrKwEGn2l
5IP2jlqOvtIhTbDNVp5jpTQMwx4IejhmAFLoPyyRyXOZyqMuuKGYCnHD5Sf+E3vvOknlk/DmSUHG
cDi0SbeJy8MjQLyD0xtP+pk9nFYO1O1DvOn8/aBRmIEsfC4bJn1xiFSFoXd76ftg1bGbGpOI86J7
KmvRdDtO2L0GbRzjtXOERSfcNm+QZ6UtKmTC1JYNk1su9U49MkN2A/+9Z+7IXQOCuc9fJ1p1kFTy
ubn6Au9NEPfFGbhL5WpFlDrkHtzV4CiLx32gzJ+XVcgZ4W63/z16wz49amEJqvJOaX9BDdhoQhSB
ZUsnqec4p6JEC6Jj2YnvbBbuz9wQfgzKyjkm1nG2pBr9LLvXh2OUt94lQf/nLX77BOyX35FUBrXC
c3ft9puHCpQMcBF6kWY0gl6xQlstgSHQJwpSYDvUXMF1mYwWJJfI2CnCOnxpvfz1LwHuaArCa191
VWP1XvfakwdLkYzCB0GOgVeMrTH07EE1fp97Lr+rvMZunqp1kfkwu9cTsSzys6i/u65/0/zw0cKT
1449jszxEE5uaV2SrL8Pu9/18ipaFvr6hWO4zqLZqhdqd+zYndEqmljuRoWGmjXlUFGeMq/Bl7XL
oSo3LLsYU9eQ1Q/7IZjhu1F4uwyW88bW3QVdzXSWebCgd1fSIuHGTtSJqDVwB5+4kmsUV3Byv4Lz
X3goNeAEiLqQRacFYlkc4nDIqxeALsylhzxGo2Juu/+7flhrlzvYgv+B58MxPCrHETmp1eMbUQRS
gy3w/s+TRvE8nldMJ4vkxSHDm+ugJpQdFLeReLp+yirQfrO97SBtOPGjAdkDeMtKeLTaIV1Y4JUq
v7ntch+8wKVjAvjM3VErDe6SvXdOLOkSKarIiDswoFmkK2a2Z9x2JztGde2ZemcyWLLcO80ca9ao
Skz3Cn3eDaPhfA0OZNZRrI7FpYOdgR1iV4GeuEsr+fzLnayTTMFMpoxuuwiXXd7nEzhJCJg1Vgsa
e6nPhif8bpe/WCQN6fKmQmIpzSkYqWORjP7pS5+iV0vJ354zLDx7upJG5Ket1PranFCWnZa299rF
qSuRNBqCuATmbLkGwTKqoBUUvD6+pM+xwj54gxkZlvj5GHHPnTPx6SQBf85sDtz8c4I044ZWDrdl
paLLTdro6e9EDcmMsHndhKThDdqIeoVzASLlXs6IlLwZpvQafWfhiiJ64Q8db/+2CiLinOaK8UFq
emuOvLPIXi4NsHV27AfW53j/zvwPvnAJ3Ej5KPhqXWHaWBwcQHeCMunsy3Hh4aKO4pDuj2p/SNj7
E/zfH81vasys9kyvbOjtHyml1U8hPyu7DJIeMSX77Lwx37BGWaJOfc47zpez6VapxuYibX5JpQZn
0QlVwmHS6/8C2MxPqFP57opC/tGpakWbWIlewwjY1V/mo4jXRxmJglS1wTgb9unH8U33lcb2qM0Q
e6pusdlTBS0UtEZkoHB14hmHgsD03tQaHKGoTbJnQcSVV6z3QFnTxNCylorcAJrEJ30fUocOR1WH
MPS2cyPM0ZGY5OoiXXOg3bggZNrsrOzL3aFUEmxMEV9s2GWTn0FbVBQFq+C6DrA4rSVmE0/0DZmA
AsDcV+FZKOnbSQ75ojky5OafocsA1pbD3plBl/Q9cGeZlu9foIwS+Q3cj0vdieICSMGaoYTqTH/6
a9BfuFZ88dTlpMDcCxa2uxIYcDvpY+oy89zdLb7oRbN3DdWGIMA1fl5RIqRm08fQz5gpoZtyq0jo
GOOZ6YLhkcyJ1d7ToDHgz6NsuIzYZupY4zRdPL/uB97DPpJ+nE21NlQXRHd8BodliUXPRdg4HaDO
wHNv1OksffoRKC6flvrpmKZ+yK9zhD1lOCd86L/Yqb9vVv5Tb++IribiH3pPWyZowN7L0Tn2B91j
213ILjRj95Zv/bomKHoCgxMSpbtn0QO8PJ8rTVmUNh/1odqXE0qUBfDuigWhID7b0gPsXXRQQdnk
03i+Ll1BgqVESl59TB/F+5a1xZB31fNtvQ2m9r4s89apgYIzfrJ2yeRu5LktG57EJqf2rIJ2issy
SOzrwHd3xIz9h05j0h4xpZA7GNQ9xhLGuG+uBvbuTXG8s34Y9eQkQm75EjYK1czYc3kt0GdkhXvs
YYYYVBSGDjna/dWKt2dsPvMd3LkPXIeQhSi6J5YbI/wjBUNNwGyEzwBkBRJVAhvGNFhkn6XpqCuB
DIdGd0Z1Is+2X4vRT4f2MW8od+hNlX801LtItipGReXFEVIXxXNjiTSTcfE+be8EMHIKpH7IFGPZ
ZNbtAtpnEqB060Y/Faxhv3V+cmjGlgljySHzA/XX3Fr9x0VZEoDJJPzfmijblQKjkdG+xPmeeW+G
ZVd/2qafxu2Wb1BeNIBGU64Qo4IvLp7SHhcmeJ/3qDB01/WA3W7OM9CCZXt0XkRicf231KbE9WEM
SVssO8QHA/w6Wdzv6lQ9XAwhHdNUKMTgBiBaqWw7ZYzh7K82HLzrpa8v1wYmkNfAdN624Wo58neQ
doTurv83a+E7ST0358J+xbXdAt/dFLLmffhg1MZQKpIm4Zf7r/mxDNjCxfloZtlMORKije89tf1l
Xyo1CmeKL4kYgv0gunea30MpyNfKqlOjnkGhuSSECeEBNDV2eT2w6f7gs7SMOb7rdII23eNjFMUQ
1vSV/8Qwm8JyMHUB1LnCgQNw4hTPsdTzzyQNXzCkJNhf07sdDEj1xRLei7jx7mvypv1gJPFBNshi
WJSgXnvV/wwwi/gk1UB1oExWEpmkdWg8SZdqNI2WYvr7gdti4RGy/6Cup14Du7vr/qg+fpwefwSM
H22kloM0fjC++DkveKUYuAAIELbbp9116IlOkUqfEONcHQMNwSQaUPLPED7pboEcS44CQeqOhIjo
YCIFFCJ7KSyMwzhE1Q414T4UblOCOvCcPCKiBwPUxOyFhlODUPDtJhPLYlp8K6eafAHv0U7pMuW7
0sWDJN1OZEsrMqiP4eHW6ckN296jcJI3I5PYfXnjpcC9YmMrWBUS0Rw/xokuCOVc0Bgm8WymhmDy
rrm1yoVVXJwUkJuwDbbhzJ2piWSQpmPZWhVdSalGczb8zDECq32GvF5KpmtZ6uzMbDUDymFfc93u
nKHUtS4WN8707xyD6KesRTXw2YDLpBiUghyx/qy1PBy0XZ+eV1Hnotav2NgH6tEVL1bpx4yKQOr0
pjJJ5RtzbysbF8kyF8oGc+TyB1RbK0pbMIi7KiO62QD41nRwBxCNdE7R8owr6x9Q02UaD+1SHQaG
WNynClBNvfYLY7GU8qpwLar6SVvKxgo+XVOZtpiCspsT0wJWazEehD25L+g1bR8uI3IIyOd8F/CQ
SRl8FiYfRt8bv7g2yqyeslCyD6UFFVkZYX3nFqjcDR3i7+ow9UK8t8LFzlivZABNEahReIyWSqWi
3/oRGb8+T+7hZRqLVcW8zzsUI/qqJ5QXS465/14BYI/7SwueOXbv4oVnBe0rH2yF5pdUtm8FKga9
uhz7+00q/i0nXek8ZPz/s63Vx3C0auJm0+bqSbh/hIDXf/FsrsCBUiX+h65Ics0JPL69wFN94tb1
oiSL1X32XggIWWjbkPAHVpMPtJ8QFVxzo7e/5ycQgSbGhTdR5Unpu/AEM3Df76la4AoQWOpJg/kU
nlSge/PvTEQjvYzeDcCrkqU1HpqeMCNmazxTCWPfGURDBCUGlo3idi/n/nGqwY3W6SzxNzDJ9bX0
v1bhqFOdgghu2BPxIFLKEBI1Xbvg+Y5Qu+lTd//NnTrEFFD42L10Tm+VZoXB5CR+NGTouY/+91Da
rAHAOOz4MZ2VrU1fn7eqM/EqH5ApJqRKyWZe7KfUps1DQbp4p5GAhICuP586P55v6qSYHY7ozHUT
oXFrvI5QChjJSRQyd1lgbcCqYnNym1HBNpGEt1JkWLg/7l592I4FAHrJOhJFgbZt5uSnrFHLeDEv
ZHBTgXK1ZgEG11TQNFe1QzX+TIt05KBS1hAWvZ5LV7asTTPl6vuh0bjEavRT7qNL5tJY2H+NJCfh
KlO/NCfsdbN9gnkF1C6QhFKSSm192vEIfXXF68CJ3bmr1Nhkum1oK/jvTh6aqSEi9602TyvFRKHb
If0ACy14lGEwJDHZLlY32UooqL8P3j2zBZmQ1eXYcQ4lfXbLHA8Cxg+EGsdKlA8KWlrT2e70q7KF
mFnUKiHb3Xaz+omS2+pMdtqQ5GIUhMbXc+CM7EwRdWSLWD7qwBmfNyeYY2ZKaCH/TeCzm7Hxm7XK
4n634/4juPzKGJIYeBfUIxUfliSBL5/bpHHCNRL2XUuyt83mzarFTP4T2sIjThxY3Bqk2wBldvS8
NQAloboiKDfg4TDN2sHjHPVF5e/Afi6/ZXmR8zyL7G9PP91IUzz8h4Qhzy4Vn4rrGDGlnfLngHRo
SmIbIRvEK1oMZmhnwKskQUYZaap4I4zTGpKU6D4L2jwJ7CpwJmtvjEri6uLp1OfCZfUhNsrdmIbP
MO3Vf9tdFtmoQDzZEJolmHvpJbOajD5txmkdVNiOkik04MGsvzmEPl4rmKMLp0M2qJ4I85tiWGTR
aCQSVKWwXCd7P+Du8eZCpuG7mSGOfpbrU5xVowNzSJnGINQKgJoOGTMckOIPW8Iv9lNYYIZMID2z
BNMggKVkKWBkJwg4ukIE/pMVjST5ItSDctmJftO/qG4+VVEWDIy6avlL01MHepSugT4g580nmtYj
dnHObQFhPEIen6paMhIa/np7ZXTL01iVpqEL9hTroIV5UnT5gj+AJD0EImRxzuQgdMrqsy5m+Ozx
pB0NLQAl6C0vlOvYYyH9gHnXyH6pI6QhqNyLmP4VjpiXiLQdDZXktYaTxOAxjHctJj7Z51MhFB9H
8VhUreNhDiV6sV8ZKiQWksbxIdgWlB5zLLc+gB4yPRcsJPeGswQPkqZDmGggwEccIrgh54dJOhP/
MIwfn0/vvURn6wMXUc5kSguluUkOwI8mAqy0PMj0mtQBC7IUiGy9HbChVGuZ6J5aydzy3vcyN3mM
N6qBv6MGkaxMVQ45GeK5YsCK3Zre2Ut/5pcyeaHjlJBPK4FBiQx3aTXrdD7jiW3eMVLjhMypsXVu
7ucbJtbFBpbw4qX2bQeoGCnwls5/l2RNkJpxkZNqh4BzkPCoQsrJPFnYL7hI0T9R0ZLcwaq3Bxc0
jHtQBGjGIDdAHvfw2rwNVYcf/QmfS9zKZiLovGpb8K3RTgPymRz2Jty5imr/3uzbSsHecH20sXP9
TZ3xVkcwFseb+DieXRfw3foQOzcG3sQmh8c9SGWk2Nu8bvpl3tY8AHqNEdPmJzjQOBVoM7/b95Rw
En4Q9e0TbTxHreUSVzOzbCcj25H0+5j1YJRVEA06xFrH99sd60Ei8RBZKhOCdcuVFZ+1mQFTqmRG
O8qGalkP5CUbka5bqvMXAiIwvH5GgH3yP91BxE8gwCGFJa1S4BKXBJQNKEVYfop7+d+oD0vvn01e
awEQrdzXj5ruKgepHEuKVDdyVBlCUCHse3NIvQiIo7Sh+Q+GMcxQwq+FvVDo8O9daVsf07qjuQOV
8yE1SEwqs6ljKQPzAzn1Y6WSCotYRkT1kzu4kLB0PeMVDB3FAqSLDTuIkaR40XryAzmuXZcBty+N
XZGaZsVuk3A8dmNTY95Y6FW41Wvikw7swCue75C1dest0eanCrp1R4QZItEs4aXtNP0abcxXa5sl
I/BK8FuGPJ4RzLc1iuxmOo0ewSYj+DnCl4YKGLvXWsVMOc/dpB63+0PHnIEUXGYx1zqLIo1JwuDx
tITCNu33FE/JWo/XE5Q5QRG9pT93rTteX1NqcJ0k4lv4eogdA6UYtPnyMfkV3SNGHQsfQP46HJP5
2TZOjx5nDERpifX9DcHjCrlTRdqXsuJT3P7w+6+c05axbuiDidz51qDcgKvGFwnUshxbe7Dj0tJd
F7XIxLcIz2U3KqTKVNIsl1pkYeq7lZhOhXavrMGlD7GdlaBmqMzW7Sm+EjKqLmnLJ2j6e4S7uO/O
65PL87jDzkn/mExhgk0+ZOCFE6tpIre8C3RXdRxzLbtI546xwBgFP35qYkg+DnEgkXB9P3xGIX0m
rD/Aq1nHrf99j0FUGy5eWzNKHsbdS8RZBasfT/btZz9Viqvxrq5P6Q00iZ/dUpiHZZG6bsHXMqOV
l1cu4IRnHd3a9RQ37D4lU0kt2cZfOjyvluoCf5Bsav3BOE4DnhhDJVyn0hhfSETGbdZsfOwjFURk
4ZRP4elF1jITbRITWXJd6Wb5vCPpmVutSwocgEgBv2FFOtV2yueJxuzmcggJKP3qrSp8/ITOQQ61
j4Ct7Z7mFTxYuKaeubWgL6HwJweRbYYi7MXjDXJ3SHwGd3yS/acjjBubuq6hm3c6BdGSfiaRX2/S
8o59fuOYBmOJkk0rv3LAJksJzSfYuqNGYX6yYflLEbUscLOedORobfHRZIammMxW1cE55sBdK3qR
Ja/DCfIZZJK1GCTfGhXPMg0Y93eKuLYznn7cgOpx4YTgXo/MhQKhsYCI1eGRFG+67Cw4zJqNLPwq
tCUOyOAn8ukTXDF4V4dF189tj6A7OO3rHq5dEhA/HPHiQYcRLn5iE/fN2/o461XV3+h7AMKkR7G3
+bOlAdmRz2w+QIVtZjp/LWOLAgxcTdS+0kijZUKeJ0o8vsebVk9nDVJsSxDlInFosiEWvzBKKtat
gHsd1AawO7SKlwaUTWps2rDqiAWbKKH4s2M3jmzvuDdJOYCZ8h9CXPzzn5X418OWO3ssWZ3Z1dH6
xg8A/ZaugLbuBYlx321h+WkRoBWyz1QywmFNEEHYTFfF3UqD5UCURwAxU4HvVwFtYdwYpFX1glQR
2W5mzk0e9eOTNHlYNbKKJLSr9wvqIRri7cv663ViDMI5OWMTvi7cWxUHJjqyarcCiI3zzAKzQubZ
th+RJGFlAgVh9s73OW23TZV5Oz+CM5Kj3g6PPV7BH0Wgtykx8QtDiGdlE/q5JzF9tv6Udf+qOcSX
pgtRxBYQMjZuyR1tDgb8OzthJWIQVII/h8ckBiyEvmJ+3O3UlGAsaj15Kn3OKIR3XqA+0CKRjBwT
uPaoWttkfuhQfO4YlTesWmls6qk0gw1nXG/JvucYvmK5IIGpzZWAPJ9fAURmGklVGjFoKverhJ9S
+lGGK4akatdERYgZPOcuL8bbKI+hdGCQYbtrZiDr4V3lpdX73aY9thoGs7h9xt1tUrU3Q8f1v5hn
FCPFZBzoJrYD0HgBhjDleTGn6wMaPyseKkdt+980liI35hO8WHC0cBHz4AsRi0L/+dyVAZw3l1j6
cK1ZUIQDmyMhYYfPGGY6ji5l45pCBkiu3n02MiKK1H7GpIUm4mZmUzSN5Wpu/v/n4SrIa9OVc8W2
j61bTgfCa/qjrFiLkEiAsB+2GXqqvaTyFMiZ+aceBTj9MKchrAkhKuIzGuAK/KUVmEsRBzv5U1An
Xl/9xxtzYtDhulr6y00Vbui3xZEbwirV3gfcd+m7ql4XMCYwKNGtrnq8nVCTW/UVhzWMVcgl4NUp
u31dECH1BotPvbJ/HoBvJ41BgeFHavhCZDmx4fNBzRRikxR3ex/CXFq+tLnrJ6P1JBd5wH9D42PP
qFKceVH8tcWVDTTVeQVJACQwPSIbWKJr1qYIEwC/2jYf2GRTdcHa8J4BeFuR8iSsSFUrlj+ym26V
EGz8JXfchsNU1NsaVL/pwnvfPmyrlNLLw5+IgWna3KW+NPuwwqhvhTAF2F+AXQPh4pHhY7zXYOP2
XXg/OrW6MnoPNpI81wuDnY23yLC8yGU9pk6yF0K/hUQnL41yyrpbNQjHpFpTtJuoe/SriIxsjXIK
kLG4HWOoJbywDLIlk53//9Tc2cW0/5G03VGYY7+WBNrScSjUO+tLzx+8sIaWNqWYB9JNXseR3cvL
Zf8iFGop4UgSVhfvaQ/9JXCxAZCUnr8EQRkV0jf4B6CqjKlqh61HIcnClhmxlTdp4vG/mpTVTCZc
h92BQYTBCpYo0fM8Mzj+kSNP+qpbmqscNwCTPI0bSdfMxGV+hUllBiwhs8F1BDEI+QGCqKR6Jx7a
iJ3sCl4T4ZJw8uX44fQPdRMNWUIgH7nuGl+vcrYaInrNdQBOnhBcyZcmpdRYjdjurcpWnheSsDmZ
ZUglG1+2eUosIcTyNoTIQplQhYquC5KNJJxZl39HPufCsJqh5zYD+tQt8TxOZhmIRCtOi31Bi6eg
jMtgoWa8eWswExsoqZkaCdrXWGddRPIvlgwDb7FTCUxxM9fbvNi2cvDbTD3PWv4HDmT5rc5Ets19
uT2ip92dyV9Vjesqso65NCEQ6LX99mzUpJVZgILv5R1B1U8aBJ9sNraIOXqm5O9q5wiKNn4+4W5m
wtQcYtMdIa6iRXkSbCxTsnPTIpY9YKzyMDzT8JVL2Mk4+KYk1zZrq6eYPK61/DrDuQJDZzipK0Ca
kPdRkiILnJJVyzQXA/VJ2OrafhkAaIxaVeYaTzT6c7fQy7SazJaxJvhFmD5nHuE0/Zkv5ZWYME+t
wbXuq1c6RrDcdsqImDK+lHa+TDpgiN6zXctr2vwAhF5q8Eqy21wrRUGeE9NRQ2SzHshtd3355zEe
r+M37KIK1xTzSLUd6DccX2DuuoaefJlEnqUfwEI6CulsalTlyyOMM1Znr33dr3iRHvpw+KhJPOdi
m+LSp61i9qQEyey65muSaPjyQuqTTnhzsiAaw/oA7A94Mk3jVQ7mROBtAUmi7pIZ0M2acLSbw2uj
0m2fCSZG8tDaEOe9wBrJwQUdHClXIc8MnXAs+ij/v5Nk9YxpAdGg75k+B1+8DezFW2lzdwT9GqJU
0fsCJuRFz+zTgBivEjD1sP4mg15T0W+oPY+q2wEN6mJvC6WRSPPtqvHc6hEykZT4HvT/jeqIOvNE
GSpg7C6h363h60/eRwBKY9RPye/Lc9wkU3kzaU/em1amEAOt8hgsEMJufXdBLWgJ+zW0dwLV9q1B
DXgj9YZdGCqbtdQcrh3+nXvdeb2vseapBW19+telRKfcdThcRA7c/i7uQDtDwGZWpKIzt/oay4ZA
hCK7vvJhxOBZn4OOMg8rtLTYkLTqvaJNIXT57DSKyu8bhgdUvDhJ4bB7SyNKRSeDHOlXapUJDuQt
nU5etCWNwiem9hyul3yrKrrY4mm+hh6eAEyUlkGCnEKeKGPbIqXRRWWGJattjtz1Iu9e3GsAi0kl
bGXLmD89ykEmT7ANQLX57730ec3HdU/Zwfndfk01WKwJLDn/1aaphGjT3iqQZQyiiiMea3EM6eDc
k+g1NeUjndnkMygjn3QJA8ZLJzux11oQrqnKTiEGfoIsJ7SfrbTD0TNfPqlNv6kEkTF8PG/yS9pM
yzyQhHpgJDrFNlQEV53UKSX63W3A8NuymTZolOPPVHQiZES6R6ezG82pOa0RkvKW/0D44aXTEzJw
R8/eorKhwo4ldmR+syt0k/GODJAWWZQ+p9Y/nFLWWCcOuaOTtyvb5Si5A0EAkDkyvrtnXxsfw/FI
/+cMZijZ+x0FEuhi4lDOkNFPkIUsk5v0M46g1IGvwS6T4e7IUudB8n/9i58mnC0a0ni7YSsf1vmh
61ayk8IBaYw4Il94tAFqfZmE+9QYYmHfQV41uCIlNDfcW0JDp30iz8LpVPBkRE4jpjY2eNBIDb7M
kiK/lWDoH1+4AflmjXb1MZGAx3gwvupSkyTBEJKfpHs2HA1ORY8t12BTfCZTXJb7NaG4ay1UV/KL
7hLw8JfaEyENyx4K5L8en5jUfiokpzcr1/dGXayHw1XaET/HuJp5YlrMmCbrA9u6KrTiRwSujP53
nefIMNEsveWRQPtlrAh0OgvFz6GwMvKduupUHcr6YhcV1RCEv9323vmPwB0w/dzST9bVFjW+K50v
MWDD9n6GvuuiPnLcXRLkeQh+SsAR/NfKLjxAhXS1g3nTzFLMiofMICYRZaELu3lu5W9MLIQ1XY4t
3+XnVCV55XyRrQ66RGDIWZPmpq9nZAoDZue8eS0p7A9EWgh2ZJyPzljsGGXy403SMzml0WUrEurM
6w4/Iet8EfSFGJwJeFbSGXHCMbcq/u4UMwTUZmPYVMuqBsAoJ2n/bp7o2YHX7KC8S0Ba90/xBr4t
Nju5QTdHQK/yw9CYR/6V5tRvZuiWQIKghOQnrFnBANc7Ric6BRdZKiNLxo6L8zEdT9NH3jNraYKP
YbnTkl0v57PnxoUL5ygkC3IbA4P1/65EsyQm7gtx2WJZYAGil6Yoe6oJETTSyrYlgj49T0CQE5fV
cVmXYUYlqErKbPVwGaBYI8jYFm/9znlHU29hvzT7+0fqJbxE9OzkgljL7ZWpSCHfrf0wf9ttWAIj
NuAi818m9Urcu+NXe7ReoeQxVMbjKUtIVm3NGyrIQnlTAKbZadSjZE5lzVSb2IFW2cyjw5AbAXyo
yeQFtY6DayuzmUGzkQUW646yT1iy1F3r5TQBCySrmgFVXLs4r00VfFFKvn41nAhGFJJ/qu4s4JKO
iPIoyD5YrJbEKWCfmGdlC03eFfgcLtmS+8NFE7lSPX5Ownuz2czJu5Sm2hruAF/tuPbLXX5rBcM7
v3Ji6juCJdArMSWnpCnoss+vVmrFOHEQzqKN8XIyQhfKQHdekn3c5pZIIYomyG3N418NJt1/RiqY
K87urgNI8f24ycyAJw5NcbwVdERwUCRtZVzQmwyfoHSIaEUka7dwZPJTHxcdaYynEIgVT8PfQV1M
c9JBW2/FboAHGZr8g9O0QlElgAXfV67feQeaOHRkUEp7DxW42eXmGGtNgGttYilQDOVuLDu1ekkI
aSo6YBjbg76V/dNBICU3KeI5B6bMcoTBysNsVGpHMhH2UqKwc9ep1+5nxKHSqi6b2gkrf+tExpMw
fYo1GMcT7hrpw8xXfIwjdmS4OaX5k7S25V6ooXqiV/01BRicDpoEiqFNyUMOpPCwXvlVJks4ozuD
ftRb0Tj9r5f7gmUSFnRuqc3mtyI4UYpGuQsKkTQURZDzLBpuzsRrSjJDwyTw7ikkVptAtVJijx0z
cnV+m1zd7Dr++kQUxmF8GulMfkm3IFCCCtaZxMzAEjT/sqbSG3zRel8a+vYZWXv8RUUcbhnU99UH
oYSOw+M3bW/S/FpQreU9BtgPlY55s20gxVd16ctEM6/negz95qZ7Xnc1AYFjE1HvsKbh3djAkLXE
ah6lCLlxYWUU6ZSSZeNcMet+CtuSnkYtDDjzohaaaIPe+7dTSH0Bd5RA5kkUhviHJ/1nMr2Zk8/a
R1AXqy0XBkEHLEaAkpHpRKCLD64jpoeUCzkAx5Dtmgp8s517JFl4OFob0+oMGdYmxArGE/Cy2tp1
yTA4ZJZBdoLFcF2m/I4nQTU2FaPJ4Hr94fF9oKLFn4+vAKzUYhMtHqlrER2/KLSAyxBMugOCF+qH
D+4kz8i3ud2czdGveoQ1WZp28JmT/9WMKCahXI8FlKXsbNIhLucZBJxsJC8oz1sSzaAztRBaer7g
ggNPpkT0bgdMY8DNYiVflnhu/Zhi9wcUPYKt7UKLbI0VkINoTLNr6auTHWyGhG0aRU4jSx6tOlr0
EHFKHpvMPW3JzECM6UUY9zokMcfdN/U0excaTRiUW95BANWf5vujTek7Dio+CebgMK2O74Aa/ie8
64ZSxnoE7O7b2oMNbgaJTDiEFbFkOMPq1L7kid9+etptCiA9ACInQ/AKQd27H1z50haFIyuRVF3b
rR7QcnW1IloP03yrHx4rRuUQ5l3m2aFQN1sS5AHyXZB/tueBnfLXj0B0SKjl7SENBo1AsJsZg5oS
fqx8fl2pMKbmb26RnrgedavT4eyTvg/V+TBWBwiJ+IwQ8/5MrY9FYvO09ARSxZz1GbTKkuaHilE9
fWOoz/Bf5+GEx0lBPeDt0JB+dE8ChY0sRDvzRv7500iID4eGQGtT710DZ2Rc1C9gLYb5wWw9nk1o
KbCGtHwJTIsFkKVrhuBrdfdPfbiDwrDQMaIC837c86svkJ/4XjLaA2wCDYDQTOLd49J88uWH8wup
LSxeFUTprcZqMXv0bBS2QtgDKhpMAIobUaxJlPk0Yzz2dwxre0yf1MVhMZicTSGLbuoK7pe5WfaN
2hmzJHgbGu1Q69mrYglDXMpi0HG2ifrf3vc/ONcp0ieCw/QpCaET18OCYJlU7tdBLGcHivKc43tf
lCQ5AzY/vodBH3Bei3pvqclHetqcbwxcU8gNyX/pHth27s4uql5iRmZe/3ajZ9akvlXkWZazQa1Z
WN3AxgtVsVc/HBamKXNp49Y/sGYcJVuCPkPepqrDUvU8HPoO08ImQjmv/9z2uAIUp+Epg1t6vZSq
cLHXkgZuGQBL632QDTKWIFizdUktBf8qmUsnnOPg2xJODZyCIYjGEuWZ6VgdbI4xZDcI7mON6jmf
ti2bqXetogDT81J/NTKgJBGEjAWa1zjgu9GulBHIfc+EHaNhEtSMxH6WG/G6dLCeDG412rahCojh
9hsDcEqX3TAeQ2by2hn1ecQ9i3w8ys3xlH5x3Swaz8V1JmasGB4zsOwSW/cFIyrrvpmNtHeozvGQ
5mERq0WjZa8hHKHOGJU86WhxfnzJmhB5yURPB9qSgGWNFjiP6psi7Fx9nBc9QuQD664iv2SIEaUq
rXypa4VLInTkVUIE6fAMZGp+C5CttWYZttlPYnIbSi+x4CrxG0rux7iuF7cJcFETOGQo6hWxfBsW
J27zpQ2sNHSdi7wi+Y7QMfHiP8UWMNnVBWbddPN2UKDZqxVTADaE9OLXy/BhJAT6PEz8hqcX8KLH
OoLq2+z0bbczi75B9muC+qWG4g7AxY+Pq58B+LuuauV331/SnwBeQEPWGGJOq3ZgtqHknf1LbiF9
iJ13G1DBwN9RVKBXAh6c2FYJRLcf+OBGXidBBaY72xwTqMxS5pwYwBf0YlfQ4R2idcqka9FkbvMR
nGaKwV7lQxCMu8hq8BzeeHk6Wc/+3p5EfDQTxD6+rR8JoPd8Q01oSJeBCU/7aGjy6QQ5uIqVbYKr
qHWJr9evSJkThgJzUq84to7UukyXDNa99sNR9cKH1A+qiCStwmhFZYl88hl/p9V4/XdnECGab8VN
QN1Mp92UoP5DvG8g+alnpobSaOPpayTMrVLHux4ESYA8mJn7QhTeZVTXijSwLpE3EuWJERBXEjKL
snK6epTHDRBQPstO0VXqE0rkpbRF088ZuD1LI5f1t7QNe775nyDXqC7aeE24aaP5cbG3c+iGNZY7
j4SOeFFNtvN9VnUPch4GXo4DzYl/aAT2XAIy/+ckPDDJNac25cFQL/RtjWJoCwU3rNN91otFYAAt
TWtaa5y4ZfzvVnbxVi0iS+F/X+4aBff/0btN5ypTnvY1MOD3UObt74gYakoljdG4QCIGKnSp/uiX
IhZtPLsEG/dFVgji7OirtVDUUai9uMJG3WxgakWyDTs9+PH6K/wq+xkBlc/veyWs8BcILeDOlpaY
C9/+ngvsE9gW6lCxyJdlKQ9HhgbgUOfT6CGPnIyhR671lYewd5PfYsOypt6HFZI+i2AuMUdvA0Z6
3QhVDyByf7UmsE/yQwJ3qAH6LFX1XZXhf40fBmGgAPRemIVyC4p8TjtHujs/MrRECsxf9kXRnaYk
Ejty/1oQIIHZGOX+9Ble8VtAZziJ1j5TAy/o7klnqy8C+zsvOkCEDTnyxIkNZs+Bk070sF2NLgNG
Rf13H10/1+/PPFgCuNGY/YYguCMLk4ZRqYJnxclXhB5guf8jty1rh2TutZK56tq1thjXOBFhPFrP
tyn1esnGNvvrduWM2SXLPk6DZf4vPhQWwiHfVCYZledmUP9xxbWMH6WJhRpjXV8kUB1K7YX2MnjX
XWyYl7Z4kfceg4UEBhqWME+DOgHL5f74/zXR6xg/wcvBom5ddhV/cSy3/v5H2h2jc6agE0MOyFIW
+V+YIkg0VxGWq10HIBbiKzpyBswRn5xgYBTUpslmP8MgRZhfzo5WXcu8kGgnQAb6r/tYKOOcbyZR
yxSNEwwUm7wpRgOqhm5DfrroXV+bY3ehXeg6CI/arxJwRdWku7XA5fwkApyVZopykAAW2Mxrp8pZ
F01gxSDuMUnoP4DNZc4tZYeIX96905PrAKrUvj/CBTLe3ENM1s4sY5f/Su4kC1k3q0eBOtadDmPD
aTkp49dyO+s8m0pNdR3K27lzF2jelOWT+Pe4lJBz4vTMrhSmuU95IoHd+3ZRDYaT+wqsmufBi02h
40idCX+IfnHlIe3aUOQT/FhzcLQjKvuwKxA22303Y3niXBSjtRD8WpkMvJzAAbSkVwMcGlA9GgVj
NEGgD7vuzv6iAv0KdNCy5cqZaqpKTTNRWI8pkjhrvTJl4qhxjlqTgr6vX+W0nvIEVZdwZG+K0T2d
GA5Piu5o73NaSRtzQT93Jq4VR2G01DsRE3TKYnkE2dxi+ge9/juyXiiP9Y0gN/4Umt1UCdyryVzD
dOVakmfuZUehHiXNWA+FY16l7hIM2Td9eKQySbHOh8Jq5R1BnqeorYyDSCPTzWnQf5WZI30+qdMj
Mu3ekp7jMO39xW5DKjbIKlTF1dKlRErOVbTLkfGrnN9QwkSfkHTyJSaNI3GuylqttQ3SS2xMFxJs
4WRhqf//Y8ZQ9cQ7eG7ZXO51qdu/UKIiNHgZCte/BQboObV4ECPFOZb7HNV1+Rg6nZWlLuwAX+lc
AdueqaTgNEzT77SXTAcf5Wj5DxC5ErgAgBwI1NRfCHvLr5GPWX9+N7BFEeTdAZoC1YkgkRnhYcbQ
REZIeS9ztgVNMJYQ/oZEBHnWHhYSoNUJU2aXD0+a/nM2WQiSoM9PkeSFXFF8wRN1OwdZtg27itUm
SQfPEvpPTeR7bDlGmFDgn+q4Z7bifORoVTTEWTMKIMWQENUS6m0MnI4cRkyC3ctzp8grBfg3R2nF
bNw7AffqVNps4T5HDbnX5HedBrVoXzOVHQf4B+OSCyLXVoHm3+cQBb8vOA7daHxaWQiobwOiigUa
5ALrLRJIHq8iwX9MhFWmRUaR6iTcK3Vicw2ZuSZBJEw8Vf/LhO2xxYeVy2Xt+c0VLyzpro8HILbu
jU13ijb/v0EjicT91CdDY5AMuMJux3Ldd5egISM/Hj7sQwqPFulBXapUoczieYj7M5ismgE06kda
kohvtnDQJNT8i5qpLoZ1IM0ZdpQMWsUncAKKM/GogPxiMKg6NZAEd9KIdhfrnwrPS28LgSV0ldIW
NcK3Tq45G37zVxZ735D8Ys4u7mYoss2A+X3A4bBLgSqmCZ93fM6l2PEhJGRtBwNiPVomne+N59rz
jdSa56A8Mcq3tIjcLyB5vfjam1cb4Tin79T4unH23GzPzhwwGOd+1Zvx+z0tJonSUMIfrtWS7hk9
zEWEJkaH+IWRI0mKSGK31XkrFJ3epIsiWziFk4KQCYcmpJYD0WY0pLBFxvAbOhQopf5Mczs/5k6z
1eLD2amZUneVcV19nGaSB/LlWevADjnMMC9pcOl7ngB2ToRhFcKDFqUpNsNTNdhfPWW8SboTP7AH
lQgc5GYymYoAZrBPK6xRzJ04lmG8yIt5AspAaQqWZyyE2fuIzVdCBc9i57WyEJIWdioQbJRFXJUR
hd6AyYVQ+d4P1Ne1sC/sEIj1Wfrxloc2eYjqZIBoXTBCKqkcYal6DuzRRV5OHcV2A85pgRmi+Y5P
GIyMlvCN/0HRzI2la1q4aF6QRSH1thJC6Sw89SNj8AAcbiKz1ewAWZ2tWMAeqS/dXHcGMy61/8Yf
y28qlA4c7P7cHz2dyKP0rvXLYVETwy0Gx28fBaOKml8X5D+ioAvEwY2pE1w5+Qxa0Q9N0pazF1jq
BaqROuJ29+qjpqkwM3XD/oCGG+iH1Q/35kfuW42gxUjTwwGiAjeBpuNU+EMZQDG03Xisvz8W/IKt
gwn3btJ0pikkL/Kc3SY2NDBGeqiwZ9HYnIgjgsRgm/MaXxt9xGTiAC9eYOH4qiwHCLmQDY5pAKLO
2XTGGpFRDHPEPUeESykT1a+SgoYu/gOp8775Yu2xRIUUaNT04Df0vSud0RBu62EZyTyAFTwGYWq0
ZFDqDtndHZVctq98t3qY4W0kbaxeWdMTHL87tFXXC+5/qInbCu/Hgsc+bT0dvmiBeV/1cvySlsoQ
IKSunOAaXNtHyXsR93m0EqnoOylg+zi8R65lsXj4i6/PXS42RixLB90UaMl7rI4SQ+W+MemGz82a
kk6yS3s0xhYycL1yFj62g8Az2Mq5OTKxUUrK3eQt97F/zB3oWiKxuxukNuTYsErnaJQOfdyRSxEc
0Qth9wTBHWSsiB1lAA2GLTRllxSBvNB/uJP09i1BPSgUEQ92e9sdChwgLPQt4cB3jAOskI7Co09T
h8dZBsFLTRP3ymSecyWnavB7J1r6/prrXeeeNwDRO446KIC4UWewMB8PzwMZ0qqOcsTBsQ/608rs
z+y4yR26HDj6mgVdgszx01UJ2kRrtpmZwZELo+G7kPDHvMGU2iYNB7ZqRQ9am/MTJSUqdmHO7RYZ
4swTEiOx7yccShzfSqsJotp7cuySJ2RTrxfNMl//0UA6j6gyApUbxUwlJd8AR5fResCOx/UC10hr
bH5C9E1P8Oph2biltph18KFN2DF0Rpo8beLpJIudeFfCrK7Y3O2puCp5whLnoogyfNv1uDP38UTO
yUkg3LKdCFrgtLndC7Wpfy5LxLY3AvCtOmBFUwBne53/AssgqUoiQnVEl3on/R3xsvbiZeFCR50G
wfYReGw/+kRf5UVhzEC1BSPx9ahjuh79iNFj9A7ycHE2lunC6WhqeUL6NJYUvhL4NhU4WD7C3FcY
8T4Aya9/rgi7YuNTxljzycmBFwsontvv2QYv9xZqRqGdS9bpe37LgaCbQBasNhDFZnT9dQu3Z8XL
V658ea5ISWBvrLoheRnb5QBApl7PfXLac/hvUhOtwS46oqgwbbjUdAX0vYQIi/SCY4oLESrOYV06
l2M/45HjyYa6GMJK5MUAQAQbCf2a8V3Eim1JjL/jstZWGlFpa2i+wL686suVHelwLbbogIAM5//m
MedWwNDUuWdxufRdjc7uz1b/o7ChmvuXKFJiadQF42IyxYQU7YB6tidotdh4J/k8PFmLuyanfhdN
VbLYUOPRi7pHr2Sqm/JDRQf3EGkIQtIFgZyXeaseP5l8iBCPS5khHrJt5XH0iW7aUxERjRxD4TTC
+pzCUkPRES2dcqJInZLkTMofHhd5v7bQeQM3rL48/DCGTN3IT91LnAP40lr8yv7t+MRwiatXsKpX
nLi94a1KeaCFssViNbQfQC8Reb3SYSwJ84WuJ0GUtLvhWWhs6ACVOvdaSdWUaufLqTR7CFL5rNPf
pp3dMeoa5jb37Jh8tE0tLUzC+bZhH40InaybrLLfufMwOBrINVrOTeBWr9dA9OWtuhjYrw8zBAzp
GcGfknkC+hfyiS1XCofrJA28iNQ5X2SgfMB9HI6ZOxBZno7cBgWK57Kaxc4DAcD7cGLvIuaTEPQb
Xe6GiEAJQ7DJmaaszxPZX53X1UTN25ECcXz3rN7R9+eu3qiG1lJ4Q//GPoewvpF97IwmH11n9lTv
etBt20tWLGtoaJruC5s6RhDP12y1A9ztIDP7eAAvCtCiXwK4Ok3uCQ4JczSOEsPcSg2kWbZfiCtw
hgwn/5gMrTgqAQiVdiEnw06staxUHM64dHB1/RZUE8QpWNv6y5FcphmppJ1oz6f560UwTOZU2Gly
cQ/WNvqKUECmmUInF0IdEI9rG+CTHlwoP7bn/Htj7gjj61ORXsbacNc+pbWQkpPipliyYXkOTlKf
MFme2QJ95uZfCGy7AxqrcP0kAfyJ83HZSsGt7iwa5tbdc9VjzSGKjEWll+t2ZVR3VXzBRZgFVoSm
U/LDXYBcuxZLGpgGREPN/ved4F/XgwkyBciVqIWqd1Fk9tYULKmGYBdikEVfKUyHoipNYBTt9yYJ
oVDTRrh37bTeTRsfXVf3kXbSsrRz+l/wuxpj5jWjWu4L6NTESwkIFiVL6ra6vb3DvfE7GSTaABLD
oD3QVbvIu92oAJSjYTKbgdd/iyRF2GNMZVcEDy2PuaI1wb2zsklm7VFgLKJ2YF+ayLs++PgD5jee
b4dbyH3enIfmDJiy4rzHBq4Zj1jmx4RiOGBN2NU8FrIu6WZcTuXVJeDg2JO7y3FM8gqTXPBku2yS
nzDtxUy785bWrXdaNs0ci+wbpeCz+Uecii3JUu8mXG7q7Y3c/Kam8N0sbvhPs9C+xtl9CTdBQsRf
hyxIPlJD4lKXFm1+mJm5LzKOTjsxthaJ8wUdINYawH/UOb0m6bw4Q2hWxlf24vA7kGbu7J1poq+i
paZLUHt1rOKYFaYFjD+FOAu6OXewzl9PXZrda2OLGx64/ZsVMFWKSBW/I1LwIwLMt0cTJ8ANee51
ShyCv23i3+ml92yxl7ayxFdfJM8txUshPbNxPyddBvieb0D5ijdQz0lw6b/S9H7dVMN+M41xdObt
ze4l/cWlR0bp+mthD5X/1xNTGuhd5To5rISF1Cr1KLGifIxMpYo6xKETOCMW8nQCjjesCwXbFK3M
Yh1h/JKBBeJy73UcQat9260Rb9M72LYAR7axk2Vb05brrmp4RDqpdabRJ+xvVfu2RigNi/MXGc7n
d2W6D9CY+X/GtlwsdAwnLrmv56mNUkuB+3XIdNm0dc2NR777XztCISEUMtpnSTStBmROgLhWW3/h
rCwbYAKKka7vlaFt2GT2uz0bCS+F5X2hVLaMaNFULgdHSa7OUGB7i7fjAojganFF5x7Pl6xpxPei
96Hjg772s5M1tDFb9J966fF+UPl3XAJ+FZNYLlRL9GVX5EUA2WAHbBdaDk4FcecXb6UOQOEzlq1f
zfQbsIN3yt93pOOD+6MP2r99v8ovF8ovMzZWpR4To4BTSUjsr01e9sAsJa4hjH5GqvH16z7KVs/W
7E0WUWq5g7rJPCel2smHxj0wfNvEHfe6t+JBJIM7PEdEWdUfGZV3c5SccKAmseQszdqi21BmZBTH
PdifQftThbZtcaPqfxSELFbBH9fSYYygmSo321/zuyE3ObGAv3I/j2L0J6gMgmOEgxhEAC1qu0G2
XhKUpAYJXOfljcgaxvsCx4uD1yyxvpdQR3XbLX9BJyaeqHzNmGfMCIU9qbG3wT3+htEzm4KBPeUY
m4KQcMpwHWaLcnexdYKmnPvngX95mGsadQbMXQdzT/h7o/b6ZWU4IIxcROJpgKnxcFA+YjwToolN
5SCusYvtlNGtYm7RvWMQKpw0RjVDPcSRJ6COoTR0sgZ6nkC1DoNM+BWbofz/VdzRGKeUd7bjLgHB
r6aWCL/D3HhaB2FpIS12SIxtRaUTn6enXoHV+DDbzFJeBc13dT6s6tZXUVTDquTerKjJfFNkKCjE
Urmp7dPclGQNH0Ulhu7kR3mPx2wY1Y0RJKnGlaO+aRZ7Ny1yZePEUq9V4j1duiHzTKGTuMB/eSEq
rhYi9dSKLsi+vhgQh0zD11ZCnVeDon3i2nhyYUUGRHlLZYFtB9MJd856ESxKw2VDUmnRw8fwirp5
1okPrwE2fBB19hJ4Z7OnsunRA4V6BLwsfsFnA7C4gj3XXw9V5AgDTmO2OQhVTkgJl2qokmJFi51e
JYhG/Synzu1NWyrh4MwtBHXGw6qI9v4xlDVvU2zByYyCha6oj5XJ3lHJ9t8CYtq9qXGrOq+PmqYg
Pj/VXfVM+/+chTO2yydQqtBBNGj1L1j/5nViHqXr4JBI0aNI2gjprL0+HZ+5eXLwtWOlnmuQ1CpG
OQn+HYRpQR3SMCBVZCjWeW20aFEzeFjrn8fy9XsBIcTq4nkUUGd5MHILfEr7XiuKqMe7mBlHeCZw
zZwSgY76MjYSbuhURQcH+4yAyqa5/T+V2B9uF/tWkchsYyzfghTe2gm8ThZdFw+tavQLVJ4DmNVh
a790iZPxKTY0tfJ/63tkAGbijXTeXVCoFVw1VH6K17SQoRNwNSp8u+9YGElkFZM5lASS37E/nFf1
6ctBgqrB3bWFrmiSOEaR4d2MGRsBZAYIjK7YlWL4Mc8rPBwgtFrZb1YajqU5dsvOChAret3pH/ne
/BryiOtBCZJh6gdmpyYtTXcv7kGPFwmlJjXOCzwCkbDeyZtv0jPIfpSPE6UDP75txdR2lUK5TtrK
zON9xQNaK7SbZT3no37UOcXqle6TzgHoJKR4aQ3zw3FXEWnIqMC3llLW1PsBNrRCCNLlXXU7t5Yw
WCl6ytwIvk4mDtBTHlY7GObRefW+197mQ5nmavD/VSjELyDmj1n35t2PXtCcjU2wga13mu/jQWhl
taHilU32/zc9ojn4VdO0wjJ0Cpp4mECqWzftniK/yK3gz+XWuw2BT/mSi0xeNVRDBKJAXnQADliJ
omglyJEEPYqDVALS4Xxk2LeDQ3QCItETpHHCXcxR83AiognNjOL+wLH7UnNOtb3Pu6YiMK3RKrJ9
G5cXsg89/6ciMsUnKDs+1hqffbVMR0EHF3jmfVbM5QoKqrK3Yk8yXuY0VnvfqUnNCjpXTYBQdwmU
kT6b1k6/Xz1HKPWndGBaIPJZiK+soG0UPnPW6y2OUs1vKOIPnGCKG+R2goQviWjt6TY7j9Xopcp0
qv0IxzmgWdEyIe4QYFNgDY01mbUx0uBih2ka/HQcfEe/ASsoYWkyIamSMGUlGeEkh+zfgrgesbb6
yMVHzGw8ZQmZulqgLdfQXdYsrcRW89yTpRMu41IQqHDZfn1rR4taIk7Th/Ek1xOliiNG39pYEW5N
vIx/9y7HvZ9XKlF1g/Z5UCShruBl/FMftQaCiLZRjNKBkSvMmnnPlGBCO0+G1n2ZKsan81k3A8bv
Bc+bYdia8yDgnHkqqMZdaOyJVM4uYAF/F9Qd7EZ0/3GWNmCUcwUmKX+1igM1S3wZ4GGBw/nLRr+W
PrQ69S/nqYkRpBx3mYcU4B+KeqKDFC6O82kx+m0qv2cXAmIHtJyuzD4yD9Nprk74dneoIu+A8I1G
S/FAufuF7x8CHJZDpZTcweCEsWDX3FegpYG7VkiKJXh7AXiAYr9LSmlhHsHTVZ3RdTRjPH6yg9+q
YojMU+F2Wot6g/hT2+4RXF5SbVTcLb2CGrXUSk3/Cv45wyHi2tdNlTqKJLQiUuHG3Jw7II+4UY2y
n6RHGQeHLjXWUgcDPNGjVKuU9EGXM4NO+uvj0u57mK51+WHjH87AAwdqaIC8ARl66IRM9ZtRSIYk
ZrwupqxImcdXvhPlXoe8jWuopJ+miFq2etqY9i/L3oQo0CflMDReCyPh5OEXy//2fu37AlTwgdQX
iK4I7uRkeddDJ1MYfDHGs3CEo1CuET4+sgBRAr48ASlBPLa1aZrz7fVykVYLhmG7E0fE3tQ8Lfkk
rv3IEAjs7MeIgwbrj0K7E2aFV1no1B8FBV3vtQeDy0KkemQiY2/00PD+x10AQG+hgBriqlmIPdQb
cQsZ5HZHJz4s7FEcznchKdaiwVPzfiJYJRTOvSIiVi1APOAAZTMy0JIQw7U+qrsvRfeQwqfU06HL
Rz1uldv0lFuj5ziRixpfNaArO3A1J/+huFJOwX39BgsJulvJh1K76NubjJpMtWncGdtJo6ZjVWf1
vJM6nmNfSgnGZ1cZvMqzNt3CeL16W5TSSHjslcf/0D8/mTQyGgIxP96xmeTJL4bqTh5Ol2iVJq87
tr8mU/BzETY0KF8a6fj1OY/xlEmcMFp9FKwO7jyYXvOVFgR3jFwPzdBqcdRLcgsLuu7Y1GItUUsx
SgH5XQ7bCa1cD43ab8QdgOhwpuyP6iuHARDOunf45PH78ua+KjUOI5hcR5VYY42g9BJQAri8BzHP
JWAruhc7L8iBjljweJ2idbxAdyfMXa3tIxoDEZSB0vMQxOTDpu1ZH7u8OAm1QSkPP8zFSLINYz2X
E97IfYEKZhBdFnUw5W/phkv9oO9dC7//ZGXsNZLnd3uJ9XxiXDsQZeI2IcoTBg8X5Slh/csha1Hw
HfABwxe5FE1Fc0hWIDR4LkxqwmoUuJfGQMB6b2PT+UnTR+vRqkoKXQG4iTt3mWh5DjsFwZfyRRjr
+pu7d1E3NyYCxCXx0MlnnKpJCB14gFEHMBYHDDzNzqj2ex95Hh7ll+jEHaI829rPBCyfIDtYTeKa
+B/dnUSHEAbGIH5YhtWnkr1oTdPV5wWT7dIAojz+U53gIyAP31bDIp/Fe4Ztbdb9bXNYrFGP27PD
ymU64Yk8E0CWq9j6/Ef6D39DGLvGmqqYu+BSuBO8BvKNRO9mDN5hgZAjKVr4aCOaROr7d/31UD45
enZjxPs9cXovDEE0diW6DzLwCyk3PjSF3YaY/HUQkQY8g7ryzIRsy0BiJBnYqlOMx57TCSkzx41H
6xGm9ufOsrcYDcVeggkKIh9UATq0fofd8ZE40ZE7v3WvXwqSTBpFbdIBG8dvqWeDobtDrGA4zJIH
T9vv1scLI6J+E2Xsm5JqSbN30TyIkN8WnyyKuU9xVGDkIgaUayCrc+qGC5feeWd2I7CpUlvkfULN
Jf/aLJ1FPBoDUA38e0uYE6FAXfdmhVZfMGIhbMz3x2nBRIDuwWSzCXIHxuCMoJGNoH3c9AdYGoLq
QIwnq0/LT/clOzEVtkLvr9QucFyJDsE8XqxnuWeaYZ87+XrUegCHFd93/zWxSRcJDMOqWrjnQKll
06iIlCnuguXcQ5H8uqIjLko8BZ2DHtzMXMJacqcYZFs+AkkvaVnPZtrBp4LnAfmTZmtnMlZzgR7t
UH+qvP2U+weJWF30YsTBAQ9XxUckpY4S85Kf5luPb8CPw1Xa449nnITNFznMfNfeq09mUwXVj1pK
GhfAso4VlkEiungw5F+z4/P0e8dziw6k+bt4ObFvplxxw2T5qVr9mB6q5nquq+I5GVNtWIlRAIdr
3alZZ7Wkj/BuybJOkGDhyYzWq20f5QRPk4xgALII3zn51ZhInAS1SD1KceRTJks66NpXYvMTXB5v
1FT07xTo+UPnjGgdLMpbRr9Dq8D28KODNEI3X+JA7SVouqgsJt6FL7HeUA1+Hv6eYBu0l+ryQ0L3
4hmVJY1Iw+jCBDam1uLHJse1KEFkmxaqeXsje5on2Wh+wTOMfHW1hMBJNfEavVEp8+XSnYrcJpak
I4WdZrfrPINjb7IK+GzWzS9eWqw0ICx4tDsz9YgwydZ7hf49/oLZafqGkHFKhOa/E1szhBsReum2
KfYn7KuW+DdHHF46cUxr4OlWGyYbuBCoo6mzJ3IjY1a/iPX1TG//868WcMTVPuAtiWxpi3wBDay0
ctwPgu2Yji1wAx1B3VD4MtrcWz0rbL0XQzsHUGSj+EjW1ulJ+T/3iGLjkWTyWmAJPitp0Bk61wpr
kTLEoxkyuTnHz0w1kwjmH5xi2kJm2b6PlvDO/sddBFaNvG8l+MsQr+d0iluDn9WDV3BIxMng3bL1
EJoAt+kBCt1i2vK1k8O1woBCvKS4orLEI2u1a5aPQtfj2rBXO4w3b7ZDLW2ORMCL1tCymd5hViKs
yOhQujOeWv3BXcLI95/MDyIEigwR5ON98kdDwlyGMSlPi1ew5Q0xPEqwyXvu8VLA1pAyNUEWN7Lk
oYHK8xLEtpvjjyauQikuELC/dax4UNHfsOLO/rTx6HWETyQ9So8UDJBzA0Wefa0eKnZgvSFP3CFs
Ok518ziKzdDLjcFszUrv2TgpBBA+jVS9A2BcuxkY++VBc6oT6vuv/FALMaC0EYHlS1DOZ7piiXuR
CmUBmBuqaCQ79t9bpMrmzdChIDMEbn/V9uxInpZT56S8e48aQa+jtWYcPLYnqA31UiTh8AcGljpm
uMwrLh9hNhi7c4rjEHav3WSE9pjIhn81YuYjvjPm6YdE6FyEzB5Nomjqd5aMjWv437jUSZtOdkpQ
rauyUlaPaT0p296hQ8C80QYNxdyQX6Mt/9t37a/mmohLAu2ehzlDpEFngzMJeumbMXPtZXd1bD53
NwaYHjg6w1ef4Q8SrOsvV2YUSQ/tq0V2N8ZuVDV339S/GsAMGW18VA7/7oyCQsn2019SZhbAFswJ
4RtDHQdRJUpNnm+j16UdJ5woqGOh6JVli227BMuzQaCKOORfcjovH6WFil2+dN4RyUlFF7cqvp4G
iRBzbBbvpaYvjDwopV9elJjuFGQn1WcNBaGRJ+8G2Iq9HQDHltWcge8Wr5s/mdasDDxQbjOoIGpx
THrShcKfhQh32cmpwgZEqwWCkA2sNg5weBB5FGEQhlTc7YeUowAxYrIauaaoWoexRe7vD1ZoR2Ka
SM8czPDKOL4Ts0TA5ZKQ2KrCO4n0cQjqvAPgjPvKsAxXPlDQaJEbTa8qof2DmVOah81jReN7Vvvg
c9mUFFX8HKikJ/irARy5V/mF7zFdnJJj96En6pCwkn7uk7PlHLlP77Nf0cik0IFqPdIO99VYdJjj
uy4KUmYTcFHwLoX1HLDC0NVbnibB2uMjq6yPA1ZEl6HLVekKl/TiE5tLlc+XQsb7/S9oJHkjMD3b
9eJo8y4SkoYmFPF+b8d7m+Omy/e9cEk/aG9LOvPnerURzYaNzHv4OHYUAWWTcPP3oz04tteV1EOf
7XqqtnNRvrITuwoaQmEnmY/Am+G32wyuAuoHbM81SseMO3PuqlgI5G2P2iLApYEjbaZLxcoBKNlb
mkoexuu/IPpPdL//E5HdhYy2r9JtARCCCJcPjMQilfGL6l5okyIl5Vs/pFRowHO2vC+mhwWsTE3w
0i+XmtqPfbtUgsyIAyg7n83C+7Oxu5Fg4HaX6ixm6GPj45RQlX+PCRcJ4G2kMYbOqkiArRDKj5tT
jPkyREu2s5U2mDu0H1nDoD0U0crK4h3S5EZFzUuEfitVLL2n4zpicg9yuWEHuUQ4rd34qLQafgx1
u+9u5zTacEeTjnpgK+S75IvwtcspYk2nnrG1ytzo76xS0VogQaQZ4quZQy32YRrEAO1W6MINsbuo
PSnyk1rXRJ4njJNNzQMvFS1mKBybpe13PvUgq2j6c/EeVF0vwhLZb9/Yz9TaRgnOYuwuzi956wDA
1BBnC+6myzd1D100lAlqqWmvgkNymXee1suq76u8Ro+N5x1lu/1L0vdcL+rXItc3ygHPmigci64m
jErBcN8k1mjw6MTPHa15ByQb/W52dRakiyKYBKVaE9F/c3kQgamaxFm6Ft0Jdqx/c2UpLPT7Yx47
J9/UivIAC3TddedGnjpvM7C9ccYpyUgs6d54r7Kp1iAIBHco/6O51Ilxlze+tjjWD/YNlardEisQ
pjJOauYVMwdnCU4HbTP+lkx/JmommXJuz4xtXovZrpbYzs9T7y4oyesMOox2vuVpmx8nfz4E9Sfr
Tw8pFUwTV7IMq+MaVPPskxkHE4FvaUiokU1SSLqiEM0sxQY82ZXaB5xblEly97k8JxLZqlSXxW4u
cllpYGt9n8AlprZxiOf3khRyTKt22rP7dNIMlSXIw5tjsUFaZzIjs5a0eQRW+6j4xFRcWtVkddbL
92phjt/zi/G4FCXmaLAc+dw4IWiif8oxkRmewE0xP+7lit6LmkfFR6D/lP4bOcULBSbhPX0uS8o8
ytnAeaSOD1gMHbTWjExdK39N1aox4OYe0Kh7dHH87UzCre114U1y9Jcyj3kuJ/hzmT/AMayzjxlb
Pfmds/UaJU/aT/GU8KGx2ekjCrfeDtYiAQTdOkQ02sJ7EyJFIfdDI4hRn1hSvrXHRS0+JjG6s/lE
G3DpJZ79q4zAtSiqiI2l/tGExY/Q/ZYA3q0cAjKEGSn6c8xobhrnnG9+aEezO8+BNIfzm9EOFNOz
+wdeyncOJ/yMj1lT1XYXUuXt//1/+LVGSytMK0bnttVBOzds3EGH6nAVDe0y4dEpP+HZrTHcKx4P
u+h2hNfXebg8zn76GsDN9PvfsmAoOmz048j0eBK1nbd9rcAlC5VLn/IwEc3isk/OUGWwXdMPh2VH
Cb1V9wVAtKUiK5+pETphfD+0f0GEZaSw1FV80U5d4LE0MQjQp8ZwGqs/Ew1TJQbg1eJNhQE0GZ4I
ZT03KpSSBvTagvol9tc87rodFggpnG6JrOgVEwyT1adJNuHWKQ9Y4fmzhjakpfOIqQ2zEMjPLnA3
T9Xo9hR3zbU9GYcP/T2vKDQjGiK34/4AbC2JiKGG5dkFD2dsvLqq474y9lj60oXpda/cFUFh045M
l71EYFbaWxj40cPmUGkyhcnGEUf3wvznv7Ow/6WNlZ26/Y7dU1vDI6BwI95Q57b2CXfqdweDdBEL
1vBBox0KCjoAUoBo2KtDKCn9OZ5yhnI9cLZgqpO51VZNNnWnVV6YnbWUaYBXsXyhC07nFXR6zyjQ
I+2ZS0JHqKImz8yhTFlSDxNSfc/qP8ZigZiLBoVtokdGNdy7kBgKUj4hzLZfUnlIyabV76k9JI8z
5vxUqYeXrL3wCo1mHB8cVqE9GfOiuMty5P+ZGA1q7OyRXp33Ai0W2xiUAo+nyYqf6sbBVcPf9JZr
1JSV76ic5NtcXI4N1nluF38tuVJRH1kjQHTdoRhNL+oaEa+UKKr+0c5vqdBfUvF1glImi3DypIkH
5SR6StTVgo9vBmex2Z330tj5ldCvajV+BHK+5HnSEQbiIjwLyO997ZlfiI1spkH+hcPocz3HWHre
UvNSds8EX/DuFbt54uBpunv4l1SQex8UkzvPyLg3Y3VoYOfQGzTjdhsXImeTZ2qm62tqzrLDAlHx
Hy9dtIglvOzeM69ArtIPbRBl0y4butwcqYkAsLEGpZltNNuCX4U6XMsvK77fzbvCB8nyFZQuOFhn
rhweA3rjQWont1l5NY69yORQFVVjtit9hBzfuReysX8MzVhlzPsAnYFptw2+PqEXTXneG56L7mlN
/68yg3ZwHWi3MjXuLalkVVg+He3S/qYgltsbrvL1tLVUtrSDufMKQOIb9bXnrUUDwb/ZtGzPym5v
r55qTTyoTRsQFX/xQUh6YYLntc7kil3lkv+Fl+FLUp7nwKQvQnRkPnPoyriX1DrNGa3K90ZRfgC2
CiaSrF+X6LqNLjS9VB5wK5KOW+9UAlOHO0/7wVbE1j1qTtJIZzfk+U9HSF5b7oJCfn8WARpgDVlz
r0EAqtI+US+0Odf3ErsnX+P0WEcRdPDOj7dFtspkjN9cQJa5CXdDZ/v2umJTrqs6ZV4S9EnVf2Tm
KREdEFZwFrcoL2pt0SqymnhRqiTow2MbAewgCr/Ytjcq9vSdVCnORWy9uYq3B32z+5YTT1MGpT2E
4rYuDTBaGgBuxvIwqhIhMZRNI6wD3lb026bCAOCDzo+tOvIkGkBIjWfL09Cv6E46mmgVC8+3qEO+
ZDwoKoRdNKGaPs77JUt/2hRguWZGhJoc771LvYs1meMCqS5soxJpH8E/A6g5VC6jAFr8QAVskqL5
fVw5W0oPpecuMdid9wXEVTt4o9t9CfZWa2os5XB0Z3pARZbcMq+/6Fh2tnmxATGPMk0k2+wbfQwx
aUIlpo1qgJ7Wpq4haiw5AJ0zoEKvvICKuzzPR0/sgl+TJY1h8mDJYOY98TDfn1seOB1PKb5K/ZPA
T/p/ksGi6XWBfsTpOGdWQSH2EtocRGlwriq4CiV5UdnfVmJFS1ZEmBETPDaaI98dEjlh1kcm0Lms
qriSu/fxBKakHXLCUoJFyY/jZ7pLRMNSJVq/r6P2adB1dCGMTLLu8qRzlQoOrPK5c0QCL23Jk+sl
ch8FhYGU4UbD/iNqRElmtJGz2HgvUuBoS7VldO+YT6zKAPjyuS1Lk79ytGT0BYchL4Nvn31/tNo2
HII/vJ2/DbRuPTVV32OszfdNHO/ZK9s47bXc0QoqiBee+EvVGWELUMa+1zWXTXYaOdT56R8vbi0U
OTYpfAP98A6C1V62HNfnCem0HvjNlp8JiIXNKQGQ27mKkOvAE3TJBG2565qbFFm6L8rwan/FLSW6
lQhULsZy6sW0xFzr65nqmjDs1NVU6vFwpcKFh1XSOMDmkOXMja8N2RC45OcTm7IcEq3XROaFDyaa
/JvtDy1siIVoGmFlt4e8a69EZ9OJSx7brqHoarzoU/d0/ybhzVYJSQp26AWZ+kVlK+lFOda6Rtyv
9G8b+b74qfLHfXa30gLWV80+f7lt0rbH+27MfylczGDLkiV3S8k0/3eeiDy2Y5LeUKhNVOsGbqb9
IxWN/jMAyF4zH+UI1IpJh2kc5A5VtDfUUdd0lY0iL4kgwld5mp8UllfuC4/EsjwaeORCQsupJR2y
7wFn2EcLtxPqgx99asZvvzHhjuOWuzMRj57VKNNeYRRqteNyIU+wVg71KZhZ1LCkGAgu0g2fECMQ
ttEDi0z9MYTQDvql5cwxfjlVXwSUBs7QdXBxZ7HprLhI34a/+yl8wY9FuMhbJHqIOAq82CGe43Bk
LoytwOYJE5RMIOwUH42xNACTBd9RpBFguiAhyglPgcdKOQO+q5l2ZUeTWvGvWMCNt0UvvB7Z2Ued
WNb0kDdG+vkVRijXxfgLhmaeVGYwwBy2oBWT696q5emosyQFM2FJXJYkTNG/dI+9kT3hVEkrpP/w
mTQwte8wZFzxLzEyt9/Oh/2huwzhpy+999aoPrCl2c/e/vBUyjZimeThyJgJa/ElkzswKjY6P/19
W7nSPqXFVTglCaf3gZ1Tl5lmsIveHT6CA82o/VZu9Be5FA6Fgzorm/kAX9hM6c8EOFc8lD2o0qzQ
xgXyb7j/yKPsbFVtYJcu9ELZFMbMNjEWrDb7JboLMsulus4MB1C9D/zPI4vC00iIij78GLUdmNdV
LK/IUlRvN7PCkclIgfK3y8Ebikv6+CG3hXcFpVFdGdUZFfW5l0u1RwDLX0c28p37zzk5E7p3RgtU
beu9U3xPVLB18rOg3CGaZZvZZWCE6MfxlwcBkGkUe2bshBc/eu8jr96jvOCoDqEjXp+CH+3rGw8V
mncvEp+izHZQVY5t8b4J+geFbVmd0ir86NZhBEp6X0RBXlnBeeygfpnXIwvTTeBGvo5fllc/IEYj
TQmLFtAOPJLp5hPEhd/V+CQ3hVu459qp3XmLUIuxNVYi7vWUPnsP8/fDHdEiXLue2FIDZApDFc8l
r38U8zmFu0+CX8DFxRcs/AcxnvBCbLIzusl0eni2f5WYYHKi1rcvp1rp454MEaW6CeabrG8d00ah
9BeGimcGu6QVMH6mzIPcGMoyN8jDpz5J7PNmP6E0aciB/sHZxu5aNe1/SJ7tR8iB9pBlevuVDOLP
z//d0QpYXFSdSocEcaKyNebF1IbrVEVQhqBzJVf38Pkb4hMSDjzjbGVbPT3QObB9DhNTL1ydZAz+
ISnNO4PBSnw8PnHdHJ7udKa1JbjU79kuw8/p9uB0y5Sk8Z3LvVugaKuJCwfmPRbJ78tnm7rTQgjH
uubQDeYxoEwEd80ri/eMk0fIYXG5lG8fE6P00B+2hdstgyWAgqqs6+Gln8TDOmeMPICN2SsVh3Iy
+5wJIYz84nCQi6hzyspLcEC0UeroJR3CiJ92PxckjGUO2YreUFY7eJ6FWbz/FMtuaD9uLQCPWQ+H
VbRmwtbkNTAbb9hI7ta88nu+ioEPZbfYLuk1a6Oke926YOBCGSL7B7QfKciXr2K56IeQ8PPdRcaG
qO458e7k1Z6ZmmXimBz5DSIH9KkDX0tyVTGm1h21x0qEhgRwUgf8ZovqAn9SeWoZPKTLq25qy39M
qCrCT/qthWz5WiC6ouKpxqKbk9i9qvdk8AFL5dwy4+jXysquQI9U5TF8MEtO55wQlVqiHcXg8RGn
hfS52Z8KQ6ov+GBZN6wlpFBW+gDophzzcmrbTCUBzxPrUBCeZd5CNZ00otSe6ITTwZbJvTxgayHi
KQ4x9Hpcq4INu+q6QfpFBSVLMWbO5F7FC45cSvxTZ8sBpqfZtIveXcM1zFuwYsuPpXZL3GTa4xdf
mqbkqLb/8qZlU9dxuxIo/tmzyIGQ/zE1UqovWBOt7+p8MPHba8sEDIQNAR6AxgBkblS6kWiW954b
+ol/JI96qej+e7uP6t9Oz42ltjHvYpgtxXLBX5CAj2m12zV9adkf6B6lXrgM5rsG7So5+u5RtZWG
kZBTfVY3Gyh2UmvpsFvb7pGfzUEsuLN4Mwaqwt4csG8PikjcI7j8o/W46g6Be3e77XAPS4DJK9vd
d8fEALSVEQR7C28+IVfrDoCIBvqLb8x4FZ0kOUp3WbMSLTEeYX5T3eaoZ5CZG198PQyo3dTiGeg6
UDtzgEStOzS8NIcPWYoFgEPtIKFfzQG5DD7wVmgngy1x1wPqkrQo6amMhLe2wuEWrVA4yLqydygc
aHmSsccXPmiOKAWW9a/F1RM78jMYXTTmQkBX6n7hSZAtuXDvAcJOjTD91RbshRuWo4WZRqxr0but
9ZR4hxBotPlx7QL8ghOReRLRZ0yjK0YTAZD3yxQ8+FOFvaerrq1gA2sbxdZA6s2hjSWzrT4lq4gb
QDwEBJDsFT5YUWIEC5Y+G0DEQQhgCbcOlDCFVqTXe43YwB+E2dm/nvSYFnzGFKwQdbtvjI+DEp2q
1ak7yyWVvrs/0DJEj2vshUYpMyrOxXm7ZDd0vMFPr8OUOZSvB3lrJsK/Kh7rJlmBjmERtVURZszQ
AgaizjFLvJy/XATgjf/OCARgHcx4nYD8SxEMWKNOwnUsxh2qv6QI18TeEDSKpMsBTHEA8v+zJJS9
6h0/tDiG6ME1BfhQnafxXLZep3P482nQMo1XUTngCriwmObD0bhnq319RgvKxvvMsBfaWLCIBFSE
EHAvFe7d1Zt+ZBhH+qNLdBvOsAxN0BIfXw92jw+ntc/RZsYPcyomB0r8OKYSUwM+/dRb4VbYAEFA
CxdvHJvw3diX3AuMNfxgVcV3ANAArejvft8W66U3ixMlj5VKbm2HZm+bS2kuzEnpf21eUdjnNHh4
fVl9HcQ8MRMeBuVphWxyc/7AiWMOMuBtilNaw1Kp7hm6JEXbmZiX/wOxm+h81BrUGE4gVWuo0ETq
CI/CAE5TTpEff/7nTNtFmwXT3Qy4KGewVvso8FyVuRUERZzThOw2K3aRLHCnviv/Q+ET4omaPg4s
GpBrXBNoQOleL+K442I0TVwavteMH8Hs7h+GCRlrEx1Q0J/qPOFkGPimbU1xFNSIEngD/NrGUoc4
Ccuc3vFux5met/no1UwIYyht8z5ftPDj1qUCbuve4xkoQUgUXaSwyjWnTHHI8/Z6NpvslRRsJuoV
S6uxJSoWWEkBPcvHYd6lRBgGycMYmTxMDp32k43WV2CLjDrGwQi4z9vDdnDi4lGvBKWtnigWSsql
JfY5W1sD93SRNWcFHDzw9uc3Q42N6NRBDuvFnyYI0jXNRqyOC/d4FfKesCAN/NO1uZ05g8jVB8BE
eM6XCtxsCDmdAEvcqCtRsB/VgHI3eOBoNwnyI+pl+OOHj/ebu4hzHPoELnJ4B+Gr6LEltkCj3y2q
EqahJzdc2UfF7uqXfIZCmF28l2afyEqfp1wW09gYT3NlBiDg5bRPVLj4g1GgDEjd8+VWw8PLM9SO
O+s5C74/Vh0EfserVXOHWavo+nfKgCEFzd/NsSnkpdhnUTIgy6L48zGDG3peWnTWLwaYmCMKo9Br
2jdYYCqJtW2QzWZ44DksAW3C1WODUB269df/gha3Vrb7TLL06JDQCH+vZLVWk4dPszWoP2qc5xEJ
5MWw2tzyD+FOxyZztzWCMBcVtXdvH4L9h0uypxtvbcjrkh7/mgw1JJyv9FG2yzmCAu1CPLkIJTTn
e4/Vp33d/iODO8gfR+5jxzaKcXyH1UaG0kQyeRNavgug8di1J7rEYoIZyBd+TmgY/NPzmRQF/UdC
rux3wUs5HmsGpkEWtFancKIvE3hgyeoLhKoVtWs+5FdAZryuNnfcyeZTliGXhSaPMGtBvtfHtyTB
OSgUYLFByhxj1OOkdMt69pNv4OH7pkOQbrdsclnF8/aU+PjczuhOZSXuevgus0/lq4/F7ZNZxexO
UVpZudPc6AM6tKY4+Zaa3cA8Zh9LQVw05HQQ5Su/6CMOZ3b38lq92AulAXS1DcSXyYn5cu77tlTS
itMrLFlqUbrKsbPeU8YNUA3n2RjBnd2n6TbPEHkpFeKJFVY/+iJ4BZ6WwpoYmz8GTEo7tPspIPZK
lDuiZOUz8bZCyw5KIlXola5oGiUuv2Qgh/XAL2GTbl+oo7sRO2lJSW0rg1Xw/UR/f3G8ZYhPt3eu
JsEWuktKkVDwsZewmRUUelFqRb5zrBCYHJMTZpMdKaeaS7oF3/rvURVplRYiG8PCOLjR+UL5vQHi
gqoRZsGa7eSYmzMpMJ3E22T8IwCd5WNr5CbPAvA22oTljolTWAAt9bA+xQt4JJP7Db9xtUo7ga8j
IcrqsxTaccEcDOA9at9QXT3n0LYGdZrjNBNdP03whTb5ttr3n2yqFTKgdCz4BDHU/rSF1I91r2hn
3nirUTwxmsewecMcuNU1oey2yowEiyzXmIUB83WLXthlwL0Bl27ldhjMM/FSYhpvWD/iu0OOBNLn
xkeoTa7AvFl1v0tvYGv0WTQFKSlMP1wI9i6YarTFLc+RL7I8/a6Jc8KTHUT75XXbVoFE0Svx9jTx
JKZ6Gm1yapl8MA/obxaHi9ZiCLIvQH3kcWX+9BeL9YydjGeRn9B/VrUouMNE7nDWVLSr/SCq8shd
JMt2ZiRgmpXsJj3XGC9QlSrOJwAOUeRq8/XIWJ4SjDSVKQC/KAaCUNZiTQ5jVOjXG3fHm255MIFJ
d9cySZMjZpEMvmtnXAprE84a0bPAvAJqCepFBLIxvvXrwBYj2rflquAyH5YAtmEIiIVZumftLY/F
KHwsVLj7w+mw1ZxGryckZRajNKwkh/EkWcudZWrWtcyYy6YtOzvK7Mk+xr8B+sAMDmfcIzDrxJU/
MDNXPsrV8C+4AfZE9ukQm4dgqkoZmReUvOiqU9dFYaIgjFaBHcMGmS1QTLGJASe1+DOrXJ6YCMFU
ALcU77id0q50XiLpybSi/wbhTIcfdvs3cOaFF2aG/X+l+UbCwWLdtfu7HNgLh+0rWrxsNRXiUgHK
of7LZl9lJr6NQHA3ruwPtdryDi2LoLZ3G6zRDDrpVXNTxmlMzD9o2JRWuUHR7i0g4r60JUc9xg2B
jQ7NRqO3UdJFVUPnuXA0+nybJyJKyOZdIZx5DtvNhPN/CtHA8pIbEYK3qemTWRLpBIBWpXBvqnmh
oyClOYaGwdVK0kk6jvoZXjlDpECX/VOmVZxMSYUNLCWdRgoiISSxevvrVrLL7V0O8XWCvrfsyaRl
qc3E6P4Cc7F8bu0VzZ/lwIsxrHNL8BcrUymRJCGRnLhA/D8kIfSCF5HVqB4kaiurgKuViGnzxuZE
xUSEnzWunsP1tfuC05VdXTbIgy1AUs40aJ8sLcmAPnWAXMxm7KsC5oFoEYuV8kKmo9zeLFFj/N+A
P8d9NT6R8Qp2R5Fr6xhSDRRrI7BMDRKiIPNM1h8aWlVyap07Pjq8SRnimLQ/d6fptFJagaa4ENDh
DVCt5NcyntMT920DTanUXYUDaHpwzBpE9rxJf3jvTiv+gdi6iY+/bZb81vXVf5FeUgIvXcJheLc2
z1XSrKjzpH5uRPqD/wT131/J3Yv5agzfiHdnfMmjCVEWBgfU7U9UYQksN7Dd3VRsSX4B0I5KRIlP
TsijMDYbB+pDoJzTYrmP6TpsYGeYUH4awSlRGt5o1Nbx61cMpwqCQyYmVm34vgUvWZspfRqd456/
9MA3TG0+J284htQtmiiSXQrOfsO4jtdim5haCEE22sa4S8mcLKCBbunvL7IJ7kCMrtYGz41TNhyg
IVn4FskjKWP5YoS2FEksm3Il76TmR3075ZC6GJ15sqWr/7qnWEv5ocK8LA9f4A83ku349Dmi9hL4
0EFmJXwCrhFZSQaIUFnE2casYmzt97r1EUplgAMQpAPR+oo5c2+rZI5UzlGiPoHp74y20gbfzwgv
v1kAQ6yxsZ8/oiaZMaYR2j8Pe5O25jHh+eccxUwu/552D/HDtMj7B3OOXF9uykWZWVg1fZXbOQqT
+vWclsFUOM4jxgEYadu8OaiNqU3Rm/IQrIkcAZDrRqqmer/r1N6BCihvWfhMy6TsIPKan/fYMT9l
jFzaW9uOpBSvJWSAJrm72dfbvkAhYjg9iBzATg8yI7zSacVaLnU802Ln/hqJMObhkeI/LoQ70I1/
swE9XZ0ZfeqvmvrH7QXdOLFjJOS8enuMF/p47UX6nioAPP2IITN4ASUxR++nMLE3E5/hI9GoNBL0
t3mkkxIWrZKKXCfCc40DCXPJS4/W7jUvfpbbp/F2bMsTSxPdG3fakBb+Eob0vJ0Eg3K63hwq4jjN
dDv/Efbcvh7lcvLZnR/XFRvQPjE6bd4ev41AVnZ9ucfs8fOVATmckaazTUQs3wCCSyl6zcJ30wZd
IqNuMuZDetC9aPHl4uF3zGLiIJcvI5OpeZf1n1w8d8vusbCGzCdfu1+9DcyY4W0hLNuaPgj2HKWO
nGuTjMw4z3mg5Z4IM59e1fvLfUbdb2uK+E0oX9xKe4mZiV7SjslK85Hy6XzjLSudfnMEGH/DU3IY
4IP6WMEnHr8/QzcUVSlxU/iXJj8EV02ZPUGjleQTq/rPvLALnL9eOlHU5iA++q1BQryeCqWeD8CG
XxuEbndDn8CFHvkn8VBRQnpD4zNRCnb6cZorPgDLqi0Ycg9JSLGTGG/xNx4YjScNU2e/IWvDkYjW
LjqgdI8MXIP/+K7Eb/sCR8Gt35o5eSJZ4hSJQ+8w0DEU+nQLlF+dR0w67aBd/ohz7jPMqwadReoB
ZXulf0sqj0hw+ZFl3dyEIkHBCbykh9gpCLEJ/7c+paqdRTtNgZiigU35O0Lq5huahPuTIFKwYGOq
Y1CUznLp4l7zEgW6BjW2PGbarruPKvr9Z4BA7Y8K5xTSlbeA7VbTLsTLjf/12GAD4NO1goAFW9bW
HmSoWJ0V5UUBWL3J0+EPUnVOWVy/tUi/hN/5yWyYC9tX0+5pC/+3ZdR0lyyfjwOEjlxZnPSkpUuy
AoEfzMwhBnDSsq7gBpBI0LuQceu29fzBUwvriemKQyNy3SFLwSaTWgS2Qt++P8OZpRVY1sEFAzZa
CCkrY7flrindiQ1wKxkAQ54UwdIU4dYC2aEQBLESZqwRhlFqppZHNUDKFC/M6apOArIghMb8zaOk
o4kpAczndXfnw2qz9Ug0T7R8a5kXCd2e31qDcg031nwrl/UXOe5ZMFM85/vDX9KofPdwmpE57erA
biZVRifsbrFWFYoDxjc6EUWjc9gVz36JAYAFfsROzymg+utax1Hu22QfFdPnA2qciTJ5xdUThUUr
98H4Etqg+SS5Ro8zx7tcYR4qw3GF/CGk8NEPBrIRaR6mwtT8t30GOeZFc0D/J8r/5BPkAk+I+dcg
3a3TFAw17Y99owcMykGf2P8SFlxWbx+GWCY32Hmk5tB0+on+wxhRKXbXl19nEkU/f0MeBhIWshU9
BhrEA8omsdoaLkxfYFjYJ+QQpzXFPKhxgNRzdySKvOag5BTNOTFKroPjKXldHIvzC48OHkV3QvBn
9LTsRP4Plun4K3XfcqlfjHb5hDZdHCx2aCo+WqqEKOUDDMvwsyQRE4r80/F7ziqSzct/8ZGr70w8
9bjARF0AcT6qP8e4xngAXlKN+DMcawEyXVZ5kR+ovZW0dly831FhScYQRPMdSizesnCxee5m6SVx
uXCPJde/pP50haqVn57qZLX9I/u9oiwd/U8xn2a+ZIWTTlRGT2A0NUcXSb6j9wopw9WX98HdPIFe
u7Gkbhasr2PUrdIrdKYQKZwgNAOSHRFtRUAbhc8YDyHYoc7ebcgKd8qVtf8ZHCpU49uKbEwQpiIU
sFBalDL6FzuqUd7ON8JM9xbW4VbaaQgPvD2nn0bE8OSvhwZtkQnwRMsuhvI9Dh6Jro51nSRAqqLQ
iK0vryK4R/IPcpOFTzNrchrsPhr+LF6sVUExbg3SlrWsZ02lvJkUVnNvL8RURpxqF6XvJ1+SgaaN
d5s9e19j4n+rimjilEAvA9QwQLMCGuVV6+tcJOd8JvbtD0TlgpjEEfnRk/JziWX9pHpLzCrBF7Xk
4Gh6O3B1gVIOjC75/yTqZK+krl3u15uRf7iGRV4v3jTrRZZeJHfPMPK5h25kYAU43cd9xPPNhiyE
1qAosBNWV4VHQEzRvbxLlqw0XQ55XopTNyHOYimruImlhwBFvHCcr2aL9397jLMWrAYpjmJ/r3vx
41dIjd2aWI6uWd/IR6+qRb5Oxxgkk3ePZY87YN7sv88+BX/Uu/L29KrIIwPdgaRa6k9iqtpYSs0w
x/kK9kPtUaBAAThcGVD1AghWNHI/9nmCZoK3SjkYCq2Kpr0Kk4S5xy84LtC5Rqc6ut3oLpkYIUZN
NOE8PimcnO7+bTsSkcRZ9LFGXO6utxJXw55vX1/eeTLMyp+hqn91jjc2XPMqoaJG8VZtCycrXAnG
f7i11NqmGFsVPE8saEz6Luz3gC1iwPcy3EGfUjnCoXkkzcdW682p4B0c1YGnw3dwFDBCkire9pB5
un4pRJLBo6886UnieVZfQPjpdJhbHrANDSNe0/Cw8kksIL6p3ktFNAbAODTtdS8aGc/zuny+O8qy
PapRMt7s8wP9sIa3x5tSaT4dtlcPED3nFmvsxB0ldiDTOGfunlJSqrNYPXZ1zQOZrAa0RreAiwxQ
U+xFDAKF+z1+fTwwb0dxLu1UWoaGSE2pXFR2ilgqEm4nUsMtovN51LHA3PXbLLlmjGQp6jQ+qz+0
dugIofTZHA25yAzx9WGvULiOjHU0HNf9d8/7eV2UfLIDlFjlqm5OOGtCDXoh9y+HvG5GoJecnLno
yj0UT4JKM+atHVLnKnUY0xSMegt2l3k4aVPnW83iHQr3x171b0MURcdKkJMNF6olBNiSXP8Qn84k
82MrhFuAGPi1vK94Wx53BzSRj+Z6hiUMU2zgqo8fZH4vThQO8UBrU93AyKQmbVSiF9pNrpEAIZCp
M7YIk7xfjY2TUA/wC84rcyO07BSa+nnxdN1FfSLBt5/ia+QjgZpoKeLOx2I88wFd8NoRNyIGOWbf
agOL4YzAdLL5VbPkpPqSPXR8qvY+XIhxfB02OqWBgI47ibYrqE0gk9CUWUjq9fkbunEt7sInGc5D
vN/oAL5yshMwp3MN1nP5ld9lwq/VoTn5mTAHg/gZk28yTpr5ytwJNbr3D380hx4/f/CQdXqezsB2
yII+yJeq3DUlBkrNgtqMnmveLrD3k4XA5qVZDJljKm38/WclvVYI8Y3VkR9nxJbGVz3Rp2F35E7F
H79zKjYffQVFCYPbTOZL1sddjdDAI331AXd2xjZCIVtdxZ6ARbhoyViOip6OFkxmlMn3MxRsqU4u
RwOrx/V6E9fnAE0kqDZILhCH7cXF/bqQbYAs3sHoITE0v3y8dWwT2Ur5qdEkd7SkKzbKwcvgv3g3
NUaFirvUGSEWzTW1pLHV/HtejaQcdaRNim0Hr67bGGtsw5lR3p5m+a9v+CBdlKdt6OKCw7lyCL90
EhC4IQzgWzAgUbfo+2E19qxOX7gF538w7GYkA12oJxaiDz6kffSZXmwyqODwUXZ26nAFHzIfOcsr
7wk5fdfzyHiwTtHU1GB6siBtASzuFCD+7ICqkRAdvQ+S7W82K0duLFKDYH9asudBcyrP9isLp9KD
uBzfSS1NeD7WZkvn5h5Qr6LsiclDykW4yfvF6ep8D2wdI5ga+PVb0tv2CdtVOGjsD418oA2LZPDC
HuT7HjkkfHKL180zDgxDtGrwKQHoayGbjhNm4BOw3a+x4OLGoZFP6fGLrDV+ebd6LszBKrPlCjt/
UN3rd9RU1F3F54lXNMVSJ1DyP9WyIXGx3brJZtF2C+ETNIwEQHibb+BNTy/EijJzNqVrrxn4OnII
pM2uPSMYX2W5QNLqH6XWo7v7ZKmgT8fv6IWkypfXZXJMbyrv3EpR3jGm4oOTHTSYrhC+3/VPaOQ+
Mqwe2+If5SE5IaRUfC8pEKb1g5jKnXZfqIOaNVLk7wipaU6g4bJoQzgroIuA63YRrB4Hsq9eGuQR
sW9nC+C7pkaBcZ1F1oFJBLK6WGF5S9BahXqgX9JP8M6z3M9SOYoF7+natqXRBFt5i66TBPqPZO3X
JkFDDqInAMyhKuKeEgNzW4m5WMS5ctNMTVrCBObCkMRiEIpzb1VxghGNFU226UIrdlL1x+fOug6B
WETPYvy39jM5Rk764gRoV3kiisq0h/fsBCSeJfrbtC8/XgHGhrCVsnSnGlTAOhG3z8l6WOYhncR2
uIeKypU7w6/4NN7gfaBW7QrAab4A/1fSYYAQTv+s27SHrIk3ybQj124QGPiSSMkDs5g0IOQHe98/
avZnSAphyzMtAlwnyA7aY+rlUACBLXkfhk+JKuHAQb4oS5uvq7/a/y7PVOCTz6VXeuF128BUdBaE
i1v9HDgMx0LgIhgnqrDisHddi4wfriku46T617Yyv8s6e/qLH07NcJPN2+PzQWYdvfBikpwxIXaP
nsoT/iGskmOuACc75E4NixhySbmeeJQHpJkS5HRktWr9Tu4xgEvAGzzOucTE+19jP1hTXOR3qelU
0htq8tH68RNkYu3t9r9z/Du/HsBOuqUnOZRBdQQb+1V1HN108JLNJEr7vHsEz5ayJaL3ZumyJKzz
LLHXWv0P2mlQkQNLDA3hSWMeUeB29HOdPdGvc95dXvw8XH88L4nkE3wSC7WG+TcurhwzwWrXOLsa
7WUUqOlEhLYD9AgKF5W5mZTmF9bwg8QeToth8lIzSr5US5TCp1xugXpuuWEzJSeFnG0I8b8R6TWw
Uoc/6e3Yt2FdbLn1EjU2ck4Ijxr6wseJfPOJifXeiPZPc7pU9k16VKjSritb6GIJBe1qejVC6dSY
z3ECxMgoNCSO5+Rv0VrWVQktCdDouB/hOSjRjnbJC6/DIJpEY/oJiL2MizM3UVsUNu1kL4bsIHXu
gzrTgESaUKZCpOie5ZW1ORgChIXnplDwnWI1a1yrEW3Cbz1Olqy2UFbcT9zea2jFkERdvGUxP1UX
XQtO5fmZZygEIaEwKSmUPo0shSSNovHd8Q9XKcau4S6WMRfmHNoV5IjLH1n56jBf81NdrTATWWcS
j0kp7Xm72PSfXmUfrJjvZ76xi+oYANKVfsNIDRZ4V77IAKtdAGj3dF2bMz5Ojdq4pIjoYUIEASoH
zgCLzZcVcxbW2+ADviwDxTOOiuxx5GVxFJ3wVytB3ZILP4Bs02ebhm1QVsSuPDWx0hkRa0WGK+ya
cHhyObVvanIMMwu780woKpGErzglknmvm5hdYHx5jaaBXWYdPu3ceNf+WuGss3x8Ex7MNTTV0boE
6oKGew4lOxB/mnRYaMBFmy++a+EjwGBpmtgyB6uI8fbeASaoiNZHer2786bFCwuurqu+gRJvKwfH
70oEvpi1CQWI2mjiaeoAZoZTJHFOAMZIa3tSBF0JIqLuXlMDL0FHwZT6nJ/x3E6ymiB9gkWSkGvq
dp5BxkP2S6QSjlxheNA26pRyd3CqAkZR8XJafEjUY/o63XA5PcfAgN8Gsm8f4Yc3ePOs0mSOHfc0
pWIrWt0yhNvo+oZLndPwtirkUuKlMOdtORl5GOJdavopwKIQrP+zmr9NIxybMXsHlx6IrB5fr7zB
ov2MwJtfurnS5qtf2eAxpSRSQ8qKSaz9s1zM2AE3y3yIzS3vO0Sfhy2P7nXnb7subgXCaRotX2Z9
vKS9gCu+Q1NbUR0Clhlh8kbOb5fD0ItFwgyas/Wmeei2WdzuYEWpAIG1eHUVmss27JW38a8ZqL2B
+7KCQfgpE2GjUFCZKsjuFz+2npHF8FDrR+L2SzWOBRBklUrGqS40/WKqXb7z7lirSVVqs2wIttJ0
A34TDGUdvimVq9jO5ijFrzv3uA9Au41pHcO0XUqdOf5/8PA6RVRtzF7xvc5a7L/47KYep7p0xsQu
dQTVp8i59tNPH4ZOrEAnR4ETBYEPVP5WNukVp5uj+tccPm1APRBeKY5+Hbgx4IUudRo0dQsvAWr+
oXRZl+9y1OsNiG9E9r1PmPY1qMViLnLVwsizOFRs0idKz0npWIJmmIyfHJGfgGZZVQNULZN8aWaf
13ZGr9J5T1EaeKAjdbjzw2G0B1vmo845LjQk1O1YsszdW4WrhIUDFlgGg06YGppUiddLGG34gNFO
8z69vcgutEZsDMS31HkbHcDZ+AVq84BiiIicdz//j1UMefJWg594EBWTYE65vAtLxT5pzC7sOs5y
ByxswMxSnQF+wmj7GBOshhbg2yKt76W8sJCuYLbHHKSsqINWIK3JvwsfB+j4NtZanbGwNo/ZVKCb
9DcdBokotejk1LeSTKCpSLC+L7soyysnrHmNhaYmu7JVS3TCUGSYBJKQojVO+xGvn3hVx1Tv0KrM
FIRe6CcjKfTUjM7yXXxmlYUzSmW2n8J368AYk2G+2oAH8iT/GsZr6wLDWJ+NjbN/ByhUXLLq6VKx
nK3NIXNEBX7BoDnlPLCSm8UH+MNkFh1ZUvFaXhMHKAkf/k+zeiI3t45m5b8BZ1MBEsjHyoYPN4rw
9mVW7/Fxl6NdhMbx3a7s8jfsAjQSmJjCzz+Vqrj8NEND3pasEkolwAVybd10ouVNGgcP2kAWf8bj
w1+P3Few5z+IEMbzwoU/j+jf0bisk2qsd8QN7bia0xzmf94sqZq7deg75166kQORFxI01UNAYrGo
7xsenyhJaslKm7eWLBaDkl4XsPMfoYbyyCei0MPQ98er1kdXCHXom41ULJI8dwqBbotMZHDw7Nme
UN94pv9w27h5ut1DidvnASuUtXbhmqA9JK+E4u5ojpoq0pDs2Xiz3WoSSp+V/KYfgjQBDCKfkuWJ
nV5s6nu0Q4rUvaPY5ota+ihnTn+rZwRkGacDKEoAOAW3U9VxN/wWBeWX3vpI6mSxjv8kh0MYvCDi
2oa40G2h+o4/qTjf6X7C1sqyiZbwU32jrOEiiZn0VeB2zpxcRvd8KBgP8tyHoJXwif/ehrp4bKsq
KlqjXXpl/BEndkexwbZR6OnSOruHa40QsdLLvHKHX819IZaHPAC0u3QOEKzyo/fUAA59BjcxbFwI
9woC4xbLwjZVDeLnbCog5If7K8DAVXS2pVNVxibkLa1J8CRfHNtXGvg6Fao5FCesQlzY16ZPkMC/
2Af7QBc49gS50b9Z+dY/UejTZWO3O+kep6ichAe/pakRmSBB+5iQzMX07hZtU/DHoF/DDrsA3nTO
jqHw2518nq/bTD5DeWikGtmt7updQbTjWEDtjOAV2Evld9RMSPB04bBZU7XL6WlA1Hu2K71x90EP
UlqZVYnqJT2EkO2YJ5HbwC5rZYc8LM1kR97/dcT823gRJnM1XvHmh50SUx8Rj2lQ/spCJqYLWMcl
FZwQ/MLIPVFYl7jSgMWuVSk23uuzLIH7WW65B49ANQAXvXMG3GGQ1W10wupfgYJ9vLbYZ6SBt6qg
YTCsYxj5ZPLh/ZOnori99ODDM3XDj3Z0L9Zm7dFV112yc4kuYaUo8cDoFiHkJ35XH1PrJKaHb502
MNxiSTGx+xaZGNLJR8iGnjO5/MZCSMEkFBt9Ge9KG/GGoNvTydEx3yZFpY5rp92X8hoKzGzyjax7
Fo85ZUhJnKfQAAJ7bKH02nYpHwItVWUFmYo6GEV5bP6lcOycnwQyaSJzi9ogVS55jBbj2jfdZPUH
B6B4Dganyg/pr6bvRuMMwBzo1VjSwJnSyRGjJeYVcmhpCX5Fyn2dfPwUYlk+YVfxD9ylXD3von0M
vbG3mrzDRXhQVl/HY7DrWc0oLGyrKV7AIhNeRZb02cOQf0sK+D8ose4r7PNClFlQKKqc4yw/xxcS
D2dz/OA/tVAiK+hqhrgdFlAtvFMciff614kxXvTAtyPxITrW12buz1gaQzNiFSF5ZTLHybtcXVJo
w5S28bu9/+IfmeqobriQS+7QShmFlpsRKWsqdjUVDafjvnJhd+mIZc60OsnmmzljmugqkvQ80bmL
iXFZ8B/+Z9Yy/Y/MJ+SGxaPam42lfzUjI+KEmraAMhTD7ZF8P7RFo2JyfhLoqgz3dAJ/5QvISgzQ
rTge0Isv0VyFyPdIQ6F1FlybVf8s0cLj1xmO0gqhvksKws6z2ob7wUqhyOb2BqM0rQ1irr1ALGV5
pifiO/L9fOHeMdMorDoRwvoGAKAkTO3lsyL3rYNzMR1fA8MSXa7LreKO/idQ8UXVJcz8p3SGQ1UK
j6J1fNYsp3CefAWD6NmwJLgwu9NaqmPGPEgRwEXNP/RzJ6KaSGVaqvIH4RVKMeyCW1iFCdQHoow2
yrWfbrzzDU6t1IxEK72SFUgD3cihsvFx/E+ttStIPB523QrrDj6h0VSctB84llCZUx9lkYvLj7pp
+zhJ66zdJA1TVQkRVNjESnsGc10SJdb2Wr9aX2V70SStN7kg4YnHk8CCSb7bK1HntPgT26m/XgTz
fGjwfiSZdPjovtAo74H8P4vC4wf4KAGzrIcRXdZgR7Thmyx27zaOc3aNqd2ISPRupLKzDfsTI/AR
rQUyvYN7T+54U3GW3bvZSdJdEogxbWi//pYrDf0XPTTZpST76Jy8AbJg4Ac/t/MVnYEMPtO3jCS3
nlFWwombXwk5lzuaJvIuHRpM39PVbmHnlsKLAMgHKynKfLYg6x5/raFT7VrFHVx0hNiNcoemADpe
bDaK4cqrAM06ER7YVKa5zOKIzVLcDoZ/yvUwsn5gwgBIDhkyI2Hqt0cj72D8RbipJLKxBI9BviNn
k4inUyqiASpSCk7xP4+foZnHnxiMcYFcvQSAZIZPUDqiVpDG5kArAZGSG/gtOBSe0zUlyRnI9Qrv
a3Z9OJUgTdarUsZ5tQ7RVjiXmD7DDxq/K8Z9IEpWlOW2YeM5VYL4kU3RJ3nk0dD/T3axGU2A+SuS
FL+CflLyLT7JE2ExwF9BrefyR/hajXu+1/aFbWXWaNBUsnyrn5VCxh2q6o9NZ1pWDb55kyAn1L60
lxEAFfFjnopqIx+YtWwROvqKBvnP+epnl5PT1KtQo526wIPc4RucxH12hhjRatlcVAi9FBNKAGoE
dpuFDxjEA2/f4+kkq75KPRLGcHEr9DKuXamDptbuMdyBKZvhJgweu/IcUjK6suT5MRYpzhyOU3nN
4lKgegBJ5curHtvpfXNnmfypn+1n7lhCLrW9rKizJWGHNg4WTopfO17hudDxwxAEDyi2aFKjmYxv
2pgBOkIsQIsTdX5oEO6fpzY51Gwf0T23aTxdptM3fez1wppjIoO8Jp/aUkAKnYfxobuo1i+sI9kI
iQHOYH5rBFKyz1dCCb5AFuK3g32qkARxnVmK7Ml3XL22OZY1HvGmZ6MBB/yhFpG6Q4pXWbxst9P7
VtiWQyXjPsWDJCRJHLonqZJ9nzOJUjHgIIivvOemLLMT1AqjnAKdc34aLqBrctis/8k74MMUO2hw
nE5eleUWpK6pGXruUzrizvbdwLpT7EsZNxjNWebfzr1m2bOFEmE6ssmF4/MwxDSg7slibVcbYSbS
Ollu9j2KViGxR1YZ+8XQSDlv9nmaeSn1UAGXUWpbtf6yB/C7hAIrAPPeD4iL3uNMOGPDbVHojsw6
nAAJZKhqUfVCKTsmU0uKoOQpir8tMIPqVph4MfPKOZkeCDEiftorM02xa+vtZ4qIwtv7g8+3LkFM
Ml+9GGLp5cpv5fBYFwW4sEiDFQm9PBuQtdg598ATEdWXOXwSFScJjZ/RvJfft9IU1e43JPXSLe0f
cMee+K2it3EFaghhvy13v62IzsDFwHOtVX3g1IrwL6D/IAF90rNCqBSCilFtWZW20jxephK43rkZ
uvqypGCbpkzGGT7Xtw3xV2oxNwqxsv+rcomrsGo5HjmjZhgZ71J2RdxOTQ2ibMocExE6a1d4E8Rf
KCtEzNpSfNrR4DIhfP1J3wQRgza8s2d4iF8Q2w8JgUlhDjWQLpWgZ7RrzRvazOmgNdGP3LAILkv9
vf69zPexD3kTwvYNaSsczmc1+kx+m4ha8XDjFEyM80AquDnuIP12tUvbLf3X/A5p+OAK2iBmjXni
WQEEtSZVHiG9fN9Q564tUhdFrerr2LVDuVqAEz/HHU5M+wj/Q12cKsEKkwrLHH3itGwT9uYjVs8o
nPbPStdilQWBfZ0WHiNEH+8UjdJ2axz5Fs+tWo9B1YwL5J/2V3ym4T7mkQ2+eEvs1zyd+zJRMpjN
FITks5+qDdDiDMO0cP3hD7mALJ8ZZpPUI/Ct+rxXuDauRjLjUjvAQCe3JDe91bypvH6yUi0zDcKy
PSqDoOXM+/Qmf8gqP+B/Fvu9aR7tOMPANFCvwlqkly7ZPJRGfGS529UuDpYKuaZU4eUXOhd5cqdb
M51evUf+Zg/pKZmEt8SqypnDwm8GTfNkECH1XDCd8bZlj2maINYqKQQCXjUdeMjuDQk/AfjpGx/f
XRrhmOciUvTlvhUk0DFJhGlKCWvPjtV9PqykopNBTMeJNGssE6TkcizO8sJ5lLhq0oaVXj+JUIry
PqlHjkBcibdpy/qP//tkvH+p5zcBhroNjnu6vi8vyz7rJ76lvWhHMOZP/gtOrWENmmuXjZxvQ9Ba
SW8Bp76QjMoR6DcDCQpbnGIO2sMPwlove7evt26Gv9o7akGs83DH7O/FsL1+/+sLM3p10EwpIgGg
lZLDn9EIBI9IPOXczu6T34GmM+dYpdyaXUOCl6inPsVxVj8PopsoHc/yuRA25mG9Co/dP1Z0I/N5
hhIYYOCwLl032cnaRC3yQ6vbg0oq+NV1D2wghPc2bxHINI9+YF/51p9TeCGdXxQZ2AFhJjE8P0at
GXMaqnqs7LGhum0PRiqFUGESr6uwF00QzlNy8sq3ASsPkeMN3O4ApUBkII8cIvkNwC4EIyeMs09z
Z5+m0EYXQYHEiN8+JJAxbsVFq22gp+d6t1lJXiTzLKhb0Rey597GXa5y7+ZcX2E04InK8o4YI+rk
2uvjbdjB7v+2uWlPAsV8eWwHGnBE6wTwxNofN5FnoBeWp6JROHBxjvebXofteNPZ0cIKYbYnfQV5
M1zQEuY5uweTBxE44pvu82FoXT/yMLOFlvrQCJN84q+pp5W8fSJmDNI2K26uoJ/ledQglf6CCq/f
6GVQ1zDEDM4n/xilv2fqQ37eV89ZpbiQONXo8u8i7MpXe64YDBptMrQ0b6iJHZFyZmhMqXynTQa0
OZZG0g2OhKOJ1uJVb14M8VY9SYhqLHZsjHkK9hZ+Aaulid4UPHR4xTcNSE+YDO6pD9YkGOMrAJki
k4imI1LXB3nmzVz+O43XaoW2ctn8DgostTycW1Js2zAJWBa1QhZin1nfFQx+TNdXhF2wgf3bvLAD
m3YM8zMDLrQ6d3JDANJYlccGCBCyipZeWOHfd9Jsspexcy+2BzoTLGQGurhSO5bg/LPPrZYCR0Xb
fWUEAGvKX6rAmlPDIzTFV+PzAeQLfU8gCHWr1W0gH0puwNYCBTP3q4EiO3HH8TAmV8uE6KlH3kGt
itCXOzguapDPSBz7aqVYL+B9kLGcOpqVo0dRMSDThy3H77ZQS5ZM/P3bygCa76f20dQu5XJUbIZs
BN965O7JPD80aa8SnbNiOkFvn15FbYC60WYBAzHuOMfyaGgsEmvIUDnWNRJwHZLhcmRM5GRs83AR
mMOCX1g6OZ8VeAigsaAzZ4wIQeCRmw+saEegEZR3JOlox5MsAXmKrM+lyTGQuCBrePMUjQkI65J7
kzZz6pI0MOoKm8haTNlVrKLJy8cIldSHQIshBNahReuM7+JWYhTyorbvYJnjnlm2lmRvXN/1FO6L
ls/eeIC1DeiPt+oqHaQAL9qNAPS7jvQIH2fwGuJGvElwdQCE7mxmsUdy3rfG9IenQpc8h5N2pR4N
aqHI03mbVpZAA8FEMcqF2UhBypaDEMnm3nap5q2ZCvBM5p0OW1hnBJRN1TkbvMQypFAHHvnIqJr1
V1/M9Qak/1GaMo3J1/+0XLeOE9pEocigROxinebj/GXP61IcCZiS+Gcclmnux4c8Jfl7CFsfVvSx
Mt7cMMp1w2hEVdJ3jeWUl2Xb63BVdAxS7TFgL7f2MBPbPOm4poIVIsEARxBL4tREqRsyRyxe7IE6
PlsOrcpyiOTMlZhLreeVZxqPsuM32r7il/VbUkKrXYhdRweFhcv8EQUcga6TyvY+WbXKePZM8YWW
ydo7JYhTboDNSTZFPaCLFqWR4FyanYOha2r9pa+812DoEklZpn01raKlVgAuBTqycP/5N5hR9AP7
26+YCVQtZOwpyI59RwgD0lamyJHq5lPbyhBKET6hQS0ZN1/+7ckiMBZB0GzfD3P3x/ylX2rWr9nO
KnOeK2Qk/f9RPqGy7/JAJbndhJjYl62ZkzGtpG6b3CleZe8bd5mYmOuzhbTgI10Yp+xfOEUbomYl
qTuA3+dAFt75JZC3tcFD17awTCfOVzEIiFcj66nR6IJc+w4EUcfGXoodCtx3LKyUQx0VfQikpo/H
rIdh6hgpvLZt4pyi6XJMa5yJVBWm/AOyz9KO1uqqwWyayDyqHKWUHtvfKgSBehsfTrtZX0eEW+ey
kNaB+feXxF2yGZJVprMeIytxJQ6VlVMjc/HKOIn6OSYdtyrHuVszgTuRK1naV1ETRM71IZAKuIPS
NEwljwIiV+wRNhU+dzsVsFQHWW0LluqclPW4VkXp10//x5Gr1qyt92hmXPemIsCPzvkuANOpppoP
MQXr3LwPyud7vAckn9mr0HPQ8/5Ktt905hio2bMkS9jmAUraEU3xBJrxSNFPftQEj4J4B+RBxBeU
I005vqcuTBvxN+7pDqId/Hy/PzPo2yf24icwRN2koTyy9F0AaQKXqqVwEJidtbJMTVQRa+zGRsZD
gRFGT2cWrz0nAV3xJfykLOjAqzL8PQf3HyyWUgKQR5VLfcK1qlC1GhLKs1njIYxrp8wwKUpgrazC
0kpsEZr6Rc/kgu5vBokyLFCV9vTIX4aVuRugz5XSEmeAj4tvHZ2eJTDdQxGrXXlCLqYXPSX3I6Yp
ssuaU3rW87J+9Vh1h91lmtQ7nbU4zNnqHYv2tk3z9a8lVn03PZOdgj3hH5uNnwGxjvO8HqV0YPFz
7f6GZiWNbFBS7DL4Jof/FzLW5tQrG4a4q5yvhVy3eKDZQdhnxWEtDrnik/0PbxuX/qbpUURSq2iT
d9M1xXKwOwWYS/shkjVUJuao3U6yTxLefN7guC91qcu8zA05QfpnOGAWT62aEB+t8znfKRNyPhBM
aFQVudDPjAKEznZwXIIPT86suYkJuDoWCPBS2DjMj5CHT+b+U5GBsR3Ou6NquaukMUv/ZjMrHOlu
JlAPnByeVkuALh3uRqiwJ/mxVh74jcUBNp72ZTTMuLqxiT3u5vcrRHW2RvhFVs3Md1JD/fGgx78Z
EwphzYSXeaCYTFSkKpfeh3uLmqC1TYCXomT6YjisNNQvKKqe2PVcwMznr2u6lSTIqBMXT+vMPvEm
97bxg4XesuzOqCYd5qTKp04K74Jt9fhuhJC67/aeIgCpSmMECpCZDeZcgzQAjxgDkRer1tG+RjqB
cS1341xsvsSvNJXmn/VS0SWFB1TFL+DyQos2obhEDp7VgVpfDb0Rn3Vyn9KCbJkh3VVwMVhpVhh7
ScXozMGVu9XxBoimdboYao+EGj4Kp36XKn7jMLccq7k/3MF/WIEJxBTmU9tRin84d1qSE/A9Vxzw
u/WynZadA8zl+909YKjZubWJ/seHhFPnaOlWk+/GdnP0I5VkjZhCZX5sCWqxKzZpb2GewjBjcpDl
JgiMXfA1ESSMhDe8ukVbL1oT5lxnGeJlnGQonWT38ADcZ5NQIXcAOSE+VcfQ1G9fH5yiSczpCvB0
Bs75LQtR68plvwXuzb16ufb8TPeUh552mPlyOOJXt8Xdh1rAzCPlrE1lrl4oIWF7eSQg+2KYVDhM
q5xQIu6bi3qNQv1eG6u309fbmEUXdGmD1jLEmSJvOrXBdxtfb2olHjBSJidkIaw9uKz9QKgO2rut
KEtcJU15bcqmrfF3NYd++T6W2pvqJyChpZIJSLX6Bys4/Hcrb3FvF0MKCrU2+FAD0jhQ/wZOhnYM
YnvTO/aGmjXJw79A7trJ+uqT9pJkL5AJI2tA4QDZw+PAdeC/BRYpsHH9IYZAe6NoHYn5mSYOdduK
bWVFHfHYalbV7CCt26crO0DSV4cu+O5cKjarltXLxDQ+MJs2Lyhb7eMNSEQbjCTWLPlOC4Pb/7xE
bMemD24yXrQH2SzITHMbD7Uunvz1BuJ4yrblRNCAA3LSRsezhfK+nvMJFqXwRFv2PFn9tdsugmp0
7qbU1+cGnw0qaJ6cOVMVtpPUqW+amAp9ywGjXQZMJ8bldHvsPm2JJXkH1vkhadlmpujIbpw4LyFJ
pkmDQgouM4q2ISAGapf7ExUQlaFaEWudFSn/x8l1dsMUIAT9/fSEjJcESu7ulS18Rvv8lsvSOAo/
2i/c+TZX9C7HfRdzVovbs4WhYlcgGORayWCVPePfdvcCwjcL88RcQLS7tu4wpfsDpR97fZNKXYCA
sV187KkJ75Zc4pIbiJfcMCqrPEBp6l4cye3pguXCrAlGmHJzTmtaTSuYuugITkXym3T7mdc7NZC0
Ncka4FTEc4VBASq6cBRT7gpSliETRSiherilwEGZqJrhXeoVYwzY3AYi83IcrnGwVqpGt7yImN06
33jYXx/kHTzJw8cEfV/VRJMMJpbDoBecIPsgWRuT/L6ZiA+03AfPI+y/jKY51YUgwvDWGPLz/RNb
+jKikQva1lhnGczf9Ev8PMFeH+SJ+Ervl9pC0HK51rNyodBi4pYEQLiPNkrCa53e6rTk5N1cTj16
ipUyfgLzS2vM5hrv7ti+EC9JpHXfC7xVbzx74dBvHm+eCgoPYMEd0C2XsjVT3ILRRJXjY0hZ1cl7
r0tPkS82OBHLyWmq/v49fTmqpUdAHnAF8t5ee9Wdv0U9YLVaVUSpISL0EQtXirK/wmT1WzG6hAIb
eY26CslsRDqvZoh1tuzYGH7nR39hvxb4IB1lWpgEivL0fjQeuZOEzyPx8ng9TQgIgce7NZlKDfSa
1Ej4qBF7NKYKtSDtvBfQPThTY74TqZxQ0JHYFvhaqPQObh3e8xcGwF59VI0Gu/TblbNFo8rxoxBn
Vh+dXIA0YDxriAwMOuFshjNrgyfV4O4ImArVx5TCCf3HJRmYCiv2ioi+PARWUAO4R8xh0dpEqBzs
lVMDwEaPXrQ187ivpajtZrs7MVHc8/Nxz1iPIw2GvLsMs/Vg/QBU2U+sHv2potoBoxQ870X2YkzI
kqUE/du8v1+gEldsOHBP5T2AIQHSTe4RqaEcwdtX47K0ljqEb/95CtLVcOf/j6u8H4jd9y1I+OU7
4WuJtDoh6GnM/wMoejPl00ZsNiqo3uDl78LSQluRqOAOy3N0XK3ylZn2iB6EQA0ny3SOSiqS7flB
l4czlbqqLWwG6AKYw2WYUUoLDBz/WrvJ41TX270skXsPyenmQ6ZyhStAYDRzy9zr8ySxj6GocTNC
d/RZwAMB9D5wEOAiZOGlKu6OsEmcdN+prT6hiYsTAQGkU6Ailwdy/LlWVTMFcDJfSZhBuxsl8ZLL
FgV5G5nlka3MeMpOr7YtM8FlvP8FUG1gPPdCp5yoX0WUmnmhpUw6cBClZK6ep03ATB/tGL77H/Ig
KZAgD9o5znlzgYOrop8vLNmepp9fiSV90xCJwmFPtC7UKglkYmnfTXBexySrfS5wm7GatYd1F6bi
E1D/3aDqUaBCoG/3edknv7+PCHMpQXdmtZzp4sqfYOVbtKfrc7Qg970mQ3y2+61ZWY8NIc+mE3Xr
up/42CpsyEJ6yvvitALousnU9f6APX4s3515tOL03S9EWMALnfXCUJOxxwbOoKyWNIMmi8Di7oDZ
+cFumgMFUG8qsKhW8P8wC94SoMFaW2E7PDMFKNhpWywcGh02Voyy+UItm/ZW1E6y2WGpQYSpeVj0
x9RD4lFwe2PZKedvToRvuVr7DFz/N//mRohQvp3SNVZMo+z1mnd0/oOeRRG9FJNnsS5bF0I7Rw+l
UyBTSnK47wVZ14reavOqUxlXBu8ruqX0nqZfyYDAekHrOwGfb3FcM1PD8idG5qMaKM7WN4n7BgHU
kl7s+sTWPAT1VG5UER3oNFRKM45jG8RdCj7fOnu08XlIfmU5dlV4UflR+H7l307KCCkxqYcirEkp
FOsO7lm7gwJjvRP8n1maB33tOFi4r4mhszGUF67+lMH7QJ1RbiOXl8IIBmX1YqdT5pB6/GyLr3xI
p1hGD3hpyZomRCgvgraJSIsZWZJ/X+zdXYB3C4X/pG5rDcJKa+t3EZGnmbeK/4Xi73sMiBrRhLDA
ONLjLnyeYgV578EcXldbpwD5Hs96igwy7BMcztLoTcCKBr37JNocUwK1Vm8Y02kkTpe2CCOgBOqN
v9Zevq2NVJhFUcWUHmvoEBugQ1E7z0CKNEpYDSjrx4dwquQmFo2uFuvzl4s4H4MRlR2wOuKxECpb
LeLAjMPQQDObzVCdPL41zf42V8/MenxXhP9P47LlLoMoUPX4ROsRuEoapXkPcssehRVK4wsCFYyT
9kK7PiGGo0/YDo/EiZHWiBxcsJSeg4UGWZXbO461pKcvVrq4jbIwCdK8YyWRaJ9S30+byA7I4kN+
0e2wNzcZzNeRPeiCV5GCxv5ILBzEwNp767gTA7X0x2cRu7aKQEZmGZFjcnYiVp1caXJfSc4YdiIs
2a0eO6A+oe83ornV7YpYNeik6EhENMpsalr0+6DAxAs6xlXbq+QLuXttVBNUJQ7VSPLLRmUVWYMq
1115N7yoc0eGJOT/lP0UOfQzm+8Aavcz8z3lApAtimHQlid1Dz215tWc0soOO9NLsWeOgtLp20RP
slaNiOFpFgKksU/RBXw7oO7r9irrv1Hh3bpskDAYUIMB0uT4Z0N6+gIVBX35OJGKK1lQ3ezXDLBW
StGL0YOIfDuczccafeRuAJq0hA/UY8RPZAZVv+kW52SdBgFEtB7di+7h4DRL5A64XPcTn7DsbG25
yFINd+VLxPinRXr2zNaJMfzhZ3t5DFmoB+H/DgKbY2AF3cz41pvcGSNDwMYK+cqKMxKVz7tDiQW3
1SMfPHlkdaNhw33bet2A3Y+wgXxpvrQQTuXFTPcncQ8ZwvJEkdgoF3s09zAhCOUDTKgGhHfRH3cJ
3QR/RyGAmw8C56B5YFR4Pf5ZQsVoSNlLsS3fmzlPFxKc3BcJeipaRaH3uU7Mpm49xdi0SlungFfa
zPzvV5wupkbhZ5RIpFHxF3r/8GUB6EyNHZ8FF11qtqG18ahtJt13oYE9TzPYt3eN8L7wWejgrpsC
DRh3cDOaC/zaGdgcvTxG4QVDh628QCXVchfRybObEZxYsL2LwHkvWUiUCRex7fQhwNroFAUgjcJs
7OemP5sLUaQ2erS9KS5Npo4uidoqbOxu7DxnFWbFwO+clvXoBawNisU9xTB3Uzi8TF+6TUEf29S+
5Gpx6dbS6yhuhL2vcXkG8mFcfDF9Utd/+SAiwLqq0k/9N2UiOaO7SFV4njs/CdQD42XYtcRLcyhd
Jtam0CpbdnAkaayU0FyoUAQEvekXB54/2JOwbcxJmIPYhovjS8QottUOude3hksJua/bDubCPudy
Sz03qth8Y+uICK76kgft3fiDwiPCil/wYQa3l4VvUc7XQ6tB/YXu+kLqVytGNnVzSNDjvoBm9m4z
r2GX60fmSzGvGNHRyDEl0ishl8EA9nlGzRWKvhnDZIxvQe6naexnxEgTVqv5+HaQ9NQBNPpZtWY9
jg8AjSgQkmvrKHPhDbkHEbcFSuZj/otnpdeZbmo+11NzaWMEB8H3rTobF8odh9KkuNF7FZSlLYzp
LdhHuuuSHua/OxkbOzziGzSpHyHrXewII/1yOu0yg0PyEBifQZpkQUGOseVen/09U101CmG2Sjkl
YI1+O/1ild5nEnnpEHKAQxQV1+MnHgCE6NQKHgiPu73kiMwG/FIcJuzbIMxr1VfFYQnUDoWBJjJr
rpfXMIdKjLxVkCMk11gG2wPQgWSsepNHW2VyNWRTgaiICdJ3z8JNRhOvD4YK7kwU+BRlO7IoIYAP
nn8nzB935zjz5yB00gCZggd80pVMWCyy6YzdeFztb5TVbDvGd3bA5KQIbMdQJ9ZY0rJ2LuM2QEq0
/bCsfOUMa5n/ojHv878ifpEAyAKwqR+1q1qv9Qz+sbr5bOsiI4mj8JuxpEEeoV6HqZMf5FDHtDy3
Lud0hZ17CyZZEe6QX+zbT8oJECXZ+WR85pQHPD5PmbkV2HP3jC1EQNntPOI2vFDMc2VU9w3TtuWe
MbW72gfu+T9++AoEQHN6gM6n/txsZ3JReOgSk9z3S02icx/NlZDMnHZ9/bC6Rj3ZqCxzPWn+Mm/j
UJLhDLoqWqM5FGenbugf7+7hbYZh0msAxKIYs7qnFpaNoRq/1LvDU/bA2AWm9WrmFU43RndG/qE7
Vwe4UNaqHBmQlzQYM2FnTD4gomHoFvhHrnNMxVPcX1LGw364ZZnIX1lCocAdrCvFNXHjlhMCLnKj
zXIa4YPLctr9uM6Gh+Irg4C5HZS3VD+hneiqaJ7E8stMD5wvm0xM4CAeXDoxHlL3jqv9sn8M0tM/
jto+6cuYSBItpnlTUjzasNlUfzWKGQf+IOZKZ9uU8gDwziu8qfWRprxCPizNZrqzIm4uMho/1Yuk
Ji6S1nBxRpajohRmbMmzFobLlbXbaKJEyht8L9IFmqR3rUujl/gJKyyLwnUhEy4b8Jg1Av2DzpMK
Tg5qfLuclD+8TGxp5rhkSxq9zohVq8HfNUZ21nHuEwnzhVfuMIoowFELfWVNwIu7rjwylRDzmTxt
6Fo52jfYCt5myTpPkz0wpxFLeObWccGVcFOflPaEQpl45T7avwVB9UAEmnSXA+N44z37n7dJZ3ii
116bPfy7/B4iuw30E+JSLnni+sViL6nXxTFbtNWhOxfIfe/XF0ublDw+LAcIrZl7oVADu0ANRtws
ami8Ubteh3pmCacQ7O9kJFM7B/kFC4mzkUQc1pHOrmsaEgE8YHXTEYYziwiY+lEP+yt+N5lXovFW
SXKx7m7fFlX1PT3YxpEluFiPyrgeiUcmb8R5mv7OdcLYxQueJKHu/fzZ0K0tqMdbNaxgvn2ziMXZ
/9yyY/X/qXgGyAHKI/DGFTcECpJ1aQ5WL/rIjxIrqE0oRh59zfPi8ic0cb/kTE9KQkh8bQtBjzIO
va6w45CkvPxzVHJ7EWTvlPEahJaP9NSMauMzXXbCixhNi7SNHU3biHvgH+EA31yrzZlfk76Zffn3
V21KVRoB/XSf95qtTA0nfUbfSZOHipnKYa6mr9kmmE0D2ZmvPaJvPVT5Xkc85x1JIRtLLhVHmHCf
F0tzmS1LYv01uJVjxY6u0FW2/aME3bfYn4ttXzvrkKs0cDy0lTBfaZw/WisXw3KEh2T8INXoSCUM
6B7s70mkSWrmNBOAqg+Kcg8Oo6mIwEWukUNo4EK+bEXXfrHAxIAMu9BiezHMHWW4VZ763sxGTH2D
RTHiPjLhWw8nAetJRh6ATMLJgBQ92O0qblcDZ0DDGUArlTR84pqWZL27ijWS6P1TRnXLFpUD5hii
p/hmmUMCk/UXd7V71eUXn/Civb/nKKOWpz9yU8yc+XV5ke1OGWY7929hb8ErIhOmVvtT//39u4gK
/3ZYKwohg9bT0lBqnWlpBG57BlgYIoBkuUQx/j43kYuJk1tD/JpnllHmMK2mAhP9eqLXhCG1ldmI
wd27/2RWqQDcrBWnHdILNmjDApHOq4KRKjFkgVVXMjYp39qJ460L5zhuiOw9tvu9kB9dCG/oa/Aj
lMbbkUSxaEREyEfNYmImahhrCS2cImOWBrapbxvnsp0IoF9V0w6oXPx8nKXvOK+8qowD+UHomdkD
oER2oiKcx9zB8kW72bqBFOalWgN9vBoT7mziQ4J9mBOYbXjFS5Tq0duu03dnjtd2kiN22ICOR5C0
H73y9ENDpZUeDR1+eMxsM9vk9c/qA70OzzwjL4vRNrcckCrXjKlQnWleKJGUUrTuaya97P7h4dvt
dtizjVr7Y3+w8Ajskr3fp3LEXyxAirkg0BFFEfjtb8JoZvpTXnp+FFXbfDpoFDdYIuYQjUFcIgFE
t/k6GBMazIQKlzx1jwPgXOLQAXUMEjSt9vBdfht6QBXbeBuwr8PNlMX6HFTOqHlADKlkg5al6vLD
PODdBiItmBlMJhFBJPBnYp2bcX1vandmU4vQ/XydoMhymZ1aDOMHo9ZRDzwPaxvjerJZNt49dPSJ
YQgsPHVVqihqPz1xF7oXCUBTLoq8m5PVQritur0rqHbvrrSUKjSq0SQRUE04KdbS1g88BE5TcfUS
yV+QHQOtN2KVS5LwASjROJOXFvVbXMq91VCyTPEWYnVR4CcFuzH0qiPTlDk1LvcQP0Gf4ZapCi3T
PQ+MAbgakF7otSBCFXgGFSGe5RBovmfRR83/GxkcDIM5DigeyxJl87JvsHztiSfc/+s+X/7nI/m9
kDw24ufLnujOmsxho1ePzcc8Ev5ABeYPg0st69zEzoO95KQy+a5iJ/7om8mHdMQX/uJW+K4bPowC
a5qeUh0iPMDHTC/XIdA8XOp7gV8yDDPym7O5LnYp6oF1wxyiIszDl2QLVZjJushAGXoRT7kqyMdg
qR9KylXoFcA0Zahp8L0MJNpx0AMIYMF4cfpvQX2sSR28vzgBGr6v3VEcyOszhGMiyQZlX8Zt6YB0
xOGQTu45/VcHNgd/mZGkd8iCIWY/CWJyljEjBbGwvuhqsaSerkEnxfvHnv/kiBJ0fTsiR4a0XFnV
IXi3Gai9GG4NAVRIIaYw3VjOBXqQZfR98D/zJVdaPcaAE6DPB3aOkQ+PiFheeALj/64BNpNjRf7D
bRAA03X1Ui0wbrpbM0DY9QJ/TWuuOZ3Kft/rJb3+JmOSk8YAA7ov3lM5fqaN4wUK3+thtHo5jKBG
11FxUZLuCYBnNTrZOX7k7/68bb/Ir1j2X81UE3iIR1Jvz+b/0w7CFhRds3dngBI/R2otQ+YyGRKA
hlcwsEgSPgUmXWetXd6ADUF2H9aMrob9r2ctG3JrDRIle+rYY6Gc6vqU4poLR9fKlCdV60YVtpAi
Ff3OYW0K8wMSAfPWYDeFMN+6ccsOaehqdkt70LSHYYiNbA+/BdP+SL32PH56EakOpCQMSBHRswws
ZsoMU9exJtnW/f44PfJUFKKZm/B/Ng2dg+5sJwYFGKrDf22QsBYi/bnbwBm1ylzDEGoqG5TQmDDi
0OxcBrtOzCCCNcrPfqEfiaxhRlkWpjcC8+q6gjn3HIzszobneJ91OJgI2EzDIpXF2EIR3BhL8YFp
8sycm4IiJw4VsDcgqYpqijSkVPQ6vE4Y4veZtRBwSvZ2UhDCZXSzPCsBZM0UYmPajXv0pLNQjLNl
Xmm3qmq9Pv6oSo2utP505XbIrLAIUfLMXk6gM4ZIYRJcRMgurSbdG2E03ACJqoQ/GX/SCDKZrpxa
S8D6FMvtrucGnoGS6m6yIGsEKj2Gg1dDmQcRJMGENWM2sjlHKvT8OWwUruEneJeUK4kkvQvbAtVV
cTSeZ/4vFGDFUdVZSMUP8DVfTkRbFU8E20XZ8kVoLc8yoCZ8imq4Ky3E4PVSvViy57aylzOwQJaG
1st7SATYfONwygg/VyaoQvAM9t8n7HfAS+va8BAUxQ7LA2U3JbxY2f30vAsWuhInyCuqi5g/t8cD
OZzzqEQXUr6zmkgGiex3rUP4sRfWn7h6bzE4Swbsqo3ZQpenLNTJSA0cxgxo4XxJ7CcK9uMTKeM2
F+D7jk3WIYUBIgCzE4edVTWFxN7sOAm6GZKy0oqjY/J6uhnQtogFsGdZiZPMp8D7NKGfKS1fOzVr
0dbPfiJrl4Iu7bef5Or+9rMe5FVX3KK4sZPhoJAAreMU7wvVHm+Ss3qqG0h3OF453svVibIcKYZm
Zh25bVS8FzWpNOFik0e/QZ+nfkYN8dEZ1qlmoo2cljsZHXDIkWWbJcLL0c0kjdqb8VEgcRSZuzrU
wCWxB7CscSjJiroycRG2r7Ga6aUb582djj2tD2G7DjPVSdGq588SbHWsa37ag4LeQOp1J8hoI/ln
zyJvsdny2vAZYCc6Zua69Q29bIUNtGXqXks0sCLqVlIloDlJbtMugt/s9gBJI69TSsINb3JLrUw8
/Gs79MW0SiBJwFybTr245ck71xO71ZZY62zKXr/KhV/RzGLaPVY5yYQA0idiOcSZwNcbFEg11gvP
HqjHQn1IT6jzOCXoUVg6pq6jmAOgqdvx1qPSxkE0aXvioi1tmU1NpAYlWCgch5wDNywkBZqzkQ1X
n2b0mvdDmxsPg0OROuzzwJuylLKuc1XxTTwqbguumn9X3/HBDO0ZzgkwwOMx37IEIuDmBoGVm24q
aOQRl/ENrolZRutZzdSInhEGmm+7sbHuBoAJ3E62Hx53ni5+FDyCyJO/3qtICJZxipM1T39/tsdN
B1umtQZJzSb8h//hdXFT7ZhxFDXe1RTOoNfzSWS7LK/mhVwOECtgaGicmqdaJjrAmqUhLOlL0QzE
qZF3f803kpWe7hZJbOrrgGfTVF1wCa+3/i1Qlz4pEAYsMKhGmM9xEeRWO8jUK5ErZJ2Y2KN7Fy9/
8O22z1h/wYTFhpV2xyBwr/FaChA506c/X3DmKdkDsciq78dUo7FgIupcRgWLKnjsi+BHHm3NmQoD
c40awYUMVVy6rUTjjQeSEBkHQR7lIj3ukKw1d+82SIUTZI7LXGDe1F/PNrWaan3e1Y5e5LUtUfxM
lYXHyIuTXluWjlnbJ8ctW/UHpmVFWRgH7sfQ8OQX5kPWF5s+JvdLE72aG8g+JRZRMN7wfRvcQweo
DjMzxYbc7nFZG0gP97qD4U84xhCiP5Relc2VOmypvQJMzq29W/vc4LNlvgPGIQEgMgt8IwcMr88Q
XW/m4N1nEXz6U25Fdr+PRudd+X+N5oJ/+dY990/mcP8mdaErhdGXGx4LyGKNLTwm8S8gQGyMNpyr
wa3n2ZheqLfSCB6diUPJQtH0DfjYz93rag6YbwciN+afqV0Fyg5OMO2c5+plJSelZPniutQotaKH
sznW5DbjXEE7z+IvdgLZXILWlC72r5peOH0U4E3e9lwvcvXKAw9lNcEdPBgv+3swn6h0s/ai5nEL
spb2N2Tslc/f4IN66OpwRMULhouTGzyx//WKM9/mHebVM758ylHRNFo8JQp4ypdfK1kT4+NCdwvd
IarVG1Q7+eBgEewQPSC1Yz/9/kzuAUu75kW+AnbVL0w00laB3+ummVVOHxxg36MCDsiYREfdZ0Em
GDUO/9oGF1Kak7hAHOA1YaAP0acJ9J0SKYcuzbZgUorrZ4J3wEWfVe1DiMmxMactamiREKtx1LY8
UZajfOaTvtzi1ZliHvOJOUfl82XhQf43nKabPEhi5D7GgIxHAZA6h+ccGs1a+ysxocSn5VmF4LHx
xvm/724oVrNONEqUeZUIvrJc9yIUbKYmgBvlNwc59cqZvuo6uoGvads0vo4ZX/URK6PcO+g/Q8IV
d4v2J7G5/t4GgTT0lglb7WBxGpGJQ8sVQkK6fVpxCPTodYrP6l0zI4wg8ZPv8Iuiw7c7Z9UL4uoR
mDoFBvPXEiWMFb62pHbbdh2NYsOkTijOsfcE9BrMsPHvudXSn7h+n3dPxC+Dw5GFLFjmwR/8vARs
mKmTK4rTCYfEt9to7sLo5H1cOHfKSmuy/mvunmeYczCHp4oDz3tnU1I72zTlcBYsGH12HyD13hq7
4nExx4/UW9CmGErFj8vKejMSfufVrq5zZlZBGEvGkU4BHkcfx0nDxwBmjmRt2/JSieGboO9JsjK+
xShvpPdFZueMZjyx7ugcRX1UJm9wq2S7JrZV7Hyj6KhtmvZBC78cmg4wkEe1SdekYDHXi703K7eL
qqKAdUUU1+20rs1RctHAfg11pNwSdzStnLg6rz8xvRV/1Fk+oKsh1jKD1v9u6gMcT37C4qGc65FO
7uvaiKExvngHb6GIIOOZQfFKH5/4i0T5BiMoXW2maEXia2y0cxJxrwhgeloHJ0WDfoxngsmWPdt4
qX2fHSOzM1FXCSBTktl214xWxoljZB1SrUlycNaUmyFwZEYC/4anzbL3Otc62ob/pBQG8Nnrt61Y
5OuIiojhPq5xAHRruUsroxeuvYizirRSrQvD8+Xd8xrhFHzKGIJzfQ/PVoiwWhUdhdMxHBrtCNXU
U1mcMuR9gCg7aXcYsnN6f/ffxWteVmJCQB4AgM2SVG00RXMn4Giy+8SH7GTMy0//A5F/1Lh76Xcp
hNWeRi8hoXifejAc5Kb7Xy9vZKMkKJKaTciv+7ose9nXnwu5x71eaGhtfQ/8MzZdmaFziBwzYUWv
JZmbrCADTxyMtSDP2v0XdBlvlMotNyxyt6a90jQIdbf7JoLBhv7PjKLVobAzbeMEqoOEoeO6Ezha
ST/dg0q4mEQiRjPJ8Okz56ma5fFwFMxel7n1tNc+5SnxMIGLlfBsRXc+i6Q/D5wO7oTwLVTOgyMP
SdT44MoOw47/SFSI86O0JZtPbVGr7Ce9XofOddbAGFb+7naqj7QyBrrQPEbGFGFgk6DEy/fNLJ+H
CaFklwR2fnnjMZGQ6thazxdBXoyCnvpl5g90oQpro2PrvJbtheIx/0Tb2qr+bgpPEhtNlV6TOxGS
Z8j/Gu9f9vaWeZtDWq9ub1LqYc+mihQSqkFnNPRf8FEODCQcFANjZHZNGHLblgwbV3Dpojtk2YDS
H7s4sjrX4eq0DqyDBVraNe8B8/fYI5ACi/fPv++keBOOLaeO6LwCCsOMEelseHyytL8M1VGGbUZ4
8oflHEnyD8wRok8+9Q7KB/xf80nNIBSfi6iapMSMg1nxFbuSwPtBTIk0lI2RMuHLqK+alzSB6VTh
8baT9HFNVlnyQ8nEpjByv9vDal/6QKsTEvuY28DhcK9aPdZD04IXe8Twi5tDIWr/YY7lRUTpfEVP
Tbsbj760zCjqndF9eRDQQYfO5CuOiSAd0fRH25Spww6rbkvtbJ+LQuCmpbNtWLLVDgbuxOUsnSEo
8+MXyBq3Q8fmE1X6ePkBHBDcymPv6z+uzxTNdMh6B4jK9joEu680tTgWdh7X4KelqnTJwJnd5rjt
m0pOpgtqGrzdKl5pENm/4SsOuAKi0iW59TdPpkQ2H1bEcRuAl0Wkzl15Uw9So9ILJnxzx+IdNJ3X
M7dYQYfi96UU4aynzydHqAjjJTSqHbyHHdGY9Sf9UHKgCQ/O/176JTFB3fv1vCe6Ful2RuNB5Ptq
bYE35S4q+Tp+HK2Oul4pTHW8AD2A2xIGpgaYpjANjDDxpkz6BS94dRiV2A6u0EWmBEr0F8HjMhGt
2l53GefebvH0aSOZvz1HicpVdklinUK33kRStMXKuhnChTJZuDOoriH/dAi2RrLGMWgFpLXAXdax
qoXr1TkbbsDdlfJrL9u7AggxxXcmxmzPoNSbJDzewfqt+UH0y77MfaYa4WMAovyLcV/oezlS9hhv
lknI9YxYNO5eduCJLezq/1e4U+B0J1oKCg4Qptba+6rbdqtuh6VkUtss0eUM9uBV7TWd5vTaMTE+
JfEP9ZJPToitVkz8lAQCTVzoOwdYazZG2rn/pFSldLjpMhG3v4fQRFPPzsTgU/au+0LIfJ/HaVLK
EGp+xFiwuQXsOUIvMPRnRNRzXCsSdatt+drznTKgnbXZIj4IfJa7GKn1Kn+lbedFgh3/UTxBjg6Z
6rW3l6js0LRAwqa7i3rxcmDdH2Xiu5z0YoTrEfy55R3ktepqvYBKs6Z9hplZ3LJOI0P5yXcisqpH
nXo9q3qhW7Haz/aJ6MXRz3dHqyFdabjgeXE6ZKXsfTd0CyfSy2u2kn99voUsKNHh71X6/tLqZWsz
NbbEv0u2DzYRN9bDTb2dAbJWIdTmwEjwJid/mgYVrM9P1s1VDKNf87kF0eDjJrfvRi3gyRnUEVV0
HF6r1VkSSpGxSLkI29q8z9M3ndVEwO/HdsQst8e56c0GBmat1vv2M0+JK4L/5TW1617KPaRrQ6o1
LNrrW2t3/NFpsXkFuiYqjWKzFHxbIVIenGQBWJfg7wgrpL4PQIsB1besihl4/ggvNc4b/PFYtAA4
9u8jd2HrzaG0KqTQQ5lu45fDs7q4DSs28yNgSRd0LixBqMdKn4rFm3ls9dEHODkaAcGPJgGz2f1m
w0SwpkSt6qK4RoF8sASvpWRhIEbN5U5RZQtOx7KA9yW4YKWiNTUQWe+WZOuRcSkK0NQ59DncD4v6
3B91FYH0fnViAFASj3EbDsKfyuGKzHdO/dm+yhWO147UyMJtdspFXAZqhByFL6t+ZDOysl75Xs5p
smXozR0fKt9NYjkHYqvaqi/2vbFD+L72yXHJQdmltTtC9vh1mkzH8iYK8ZtlStFjRheadEgudhd/
DYe5DbZXZP/lTnSD8tz9cdLlkw78dALIN1AQTjLo1P2XFYTJMTmvoOrPgohJ+w4Aqb9vEOH5yZGF
i3hjikNjty9cg+xSR3tJ6T8yNKGj33Pe2/olwEvXt0xQ7tMJVbeUN/b4HCy4ppZxVnkn7O73WsGC
iBFGzEZIDAFVhc+a0IftaqoGBiHLyxQXnUqzA2X0+POZaI2AR7c/MsihY7h2KIEi0V+xhRU6+qyU
JS57Zom4vSAy71pu8Faeoaukq/8JUXZQPtJayJ1GyZc5gunO42LZ2oYDLLxNK9a2H1ktSN7kIUx3
d3ZypOpF7B75FXZTQSvGN+bQLz5t6q/GjMwcaIsvz2pCdV93aofbgT6MdLRgJMTa7nzyC3mhhO3r
r4yTUjEZUMwY6akoSUN2NTKLuzS5ELmWEQkScwCQ0mnChLYdQN/hbzIcGD/5dh7a5KnqiQFwX82W
g62TBF789cdaNS0AstdzZNU2tXCzeWhDyZR/c8I1fcd1uCTmAq7FFGNeUSrZETULN4j+lPD9auaq
AiL/v4G2jZC3YwtWTX6pdyhfbIwnooKOiwxnULsWqdTT1fYukld8OeuaUKn99F5May1WGfeRuwZh
sIWUIIZOzbfl7C7Q5yjOhyCyiFH5wJreV9gkP3e8d/mYQK3a1cYb0xfOWnY4kgue+NZLWvzLNjJh
og1Q47yOnHGRUH9f3FEfBTZUthknuDJAI0knjLxeV5jmvCn05rD50L3a47PbGpFVE3OvKSxXErDz
8zGjQkitkta6TTW0Me+WJtGZi1qhUxytVIfyzO1VN3t9MHiMF7qMys58rsXJ4xGnTaUtdcINxJNp
8o7yyr4aJMVx9WFlN9dWAAG99nK6Dofv8oigobi4pCii+4H2m+uLgqwFkO+0iE+6uECeMt7qQL92
Huk97HY/THUdjb5Z1WaPeRjfZMILHT1mVmaNidBbF+fEO4pNZDjL2wo29bJvwcv6pTTWo35DxDBw
dOaPqW+DYVQmZHQK+L+84eAaMzhQK/vRoEAbJcOYyqFhysL0kXr5JKVM9EEFwMU8Chys2IqN0dkQ
VEcpfNdQKy1gn/fRFyDZW3qYb16CbQiGn/dSyPg233D8nwDXbwpJ8znKCVfRKRC8QVCSBYSG63+5
SwSGxvd8MWNzH/wywt8LLNWYZlLs5c6vgGvZNyD9WQg8nOtOouq7qhW9dEjNQPibLlhPb/OoYVoO
YYIGqTnhcxUln4qtTHGLYoXeVVyyArMHw2gcJF7Ul4kWv7CpFZuXF6ykgoCrtjb0kzyXikVxpanL
XZO1SG70T9lgEsdLLeO4WFxOX7fmnsJnPcuSqJnRQkspnUBthyE7cp+ZB2jAHUr1GoLC4546R4Ju
Bt6M3Ta8MuOc2zx6Sye2IkNUgDoNBNb1Ln81zwFdtWBpwrauNhjlvyM/5szJ9QPzjLTYG/CYr6WU
Lf+JS5FT7pYg5DrMknxiZYsTU7nGESiprk7MD9fdTtVAejPzyozjc0Ltq/8sHSh7chGupzlROWlE
M+W4hsSXyCNZm7iqg97zHJFWr4Ad73TcpAp17oA3HfDW0T4HzUXj718njyWgvxpBDnSlEONOIWKN
LRiFu3COiK5xn1lH2PoBl07iE0QKlwbYF6r4B7TBYpZZGJKolHuZk3+/4/k/wlWHekTlRAmSG9kq
WAZ+EgVNKn+6zUEoe86vZsJ10zZahsJVuR3dK8gndnidErpa9/FgIVEvrKbsB/Nb5YQ3PLVnyboQ
fMRwYl6pfD/UVsLx7nWpy5SFdtA1xtsoZdRiO/h2PpmOy4jywd1pyJGOY3rsc5fnujTc6FBg162d
VExr93rmQ2xwGXGQorqhZzn3L9KS21J9zO3MAOj3YVH+1Y6dqG4AV9ZOaRRliQi0MTWwKJbPHZrB
rybF3qYOJPfWbOYKCfgZh/TPdivWFExX5Cuuh6tK86iu1DQZ5LMc0BNKdFfEUq3Nibx7eEQnzh9h
z3KhoRksoyVP+3DArbmT86ReeATT+ybQ/BFGmyEdRbWNS+tI+jHvwWnnHT0+wrcP+fDL/xVSxF2c
uD5KyMiGz6efm3A8R9s8Wzlfh53rAjd3n9QKhE0RMGU6mVr38YX3uJ2PQBUt1lE043lylgmcmkZP
rcM3GNUgiHR2xJ9wAb2UYLgPPE8w/WEKoFEX1dOQNj/3xtlg6EovUcSk25zBqjHvzArInePT68xU
xQCoNUuDHV6htb4UtkQtev65co59IFJS34Mz2EZNaNa2WHHxFYnudFIIoafV6HIiVkVol0v58iVK
/aXhffHtIUV6rrLeokFCHcWDZhgapbwoJqJamvWR0moaY1FmtFiKTaPTzyNnBf1I4zKqqsPfFGQs
l+3FDs/Jqzk8upAllF735DYtXmdB3yIY+8SWI/HGOBQlu1DgVEBw+UVyFTjGw/OB8fDtlaijBWIc
GW+J/O2jjSaMWoiKt1HvfMYnpI0ZwkfNb+Caoch+AobkhMx0w2mncQijbXkrbjNsj4YwupkLdlxo
+O/461lYYryjrp6OlSIcdn10XVmF0y/izaO9Cufj3P9Q+LPQ4Fs0jp/cex8CdYnAn2fGNc/L0auI
U3VR1FKFUhv8Q3QKEonqPZYjFSxy0InFhi+jLclTrMS33oiN7f2V41DCX5f2Ujvq7UtXkwMNN5I+
3Z9oayxEQrUnnzvcx6tmKGd1/0GNxFmV/QilPCj+CQ+HLti8bD8lZ6VLVkaCNPyezhXukMdQKA9Y
RBmCbe3okLHGjJC7+N15ZOaYA3iuuc6IGPMWQ1pFNCzvZMhnSIIHScfmgp6uzvSDBqmlQSDgZZ8F
A97HuEdLq8mkkL2O7ed3wx0t1A1IXWh74KPueChNKJQXhWZQChXPohcNyp2FAwNydWBgiil5Z8c9
OuWxITBKhjxtj7FHNPprp5eqCZKvnx8EbSBMn9lZ4oipRZ3ZnXMEXF3yzK9pN7zvmlNp7geJ+EL/
kUSiNzncAwh2zdXJIAi05/ub/O6jXUfw/yrTfPhGXPpKwTbKuPCoWmAqMLY1tbiL8CUEKWwrBpKQ
RqIGqC0vPIvPPr6j04nxLxJzo6gHwBQ6KUHstjuvyrh6ccEjqVu2aWN3U/HECjsrIZo7PRtj4FwX
zAkyyJBbygnoWJoJLTb80MqzFRuW8QeAL1e/w5zw0H4ZAdZVpmirC2NgN0fEE5DtNkg+yssOmmxI
t5GXOoIcbkNz6jG/X7KWAf+5JgIOnomr1FGgmu+3E9+LKgWaQ4VhtQxv2S+Juc9ZNJNRb0fz0x1e
x3V2vRhbxBSkXEnwIOM4mnFcN38PfpDA9bQMWDdRy3tqD/rEqqWwNb5/akp2/U+GyyvXWZ5ClQSt
0/pH5ksOD7D4dfywXjaDyMNzVHR3T/jigXp80TUoa7bE7t7rCdNGNp3K7H5aHAOleTEuCeXm1GyG
NpkqAlJXT+D/gMqmy2c4f3aj02p3m5ZqEFy9O7zlJ5mXFpOuglofDmlH8nBzkE+maAjSHQUYPcCq
l0nfAeTKZr2xYJwTD0IMERmcMCJCBSDiHjr+iNBPHmGEuh/OV4bjkcXbQIrczKTRtAU31n0ydVED
y1qPIG8wXH5tp9e74goJPEC6lFGsyvYv5BD0K3EUH+v/AlqMVWpjdvlQ+Bsz8+jon9ff04uA0cZi
/D+N2Iz1gSGrnnmeadetsuzy3EF++bte0GaXijY5qZBM7KietWx5WhBbqHR5suY34AeIX/2jZwIp
eXEZeppwuUnz5FbjoQdlNd4Edpvrn7IaHl606Lgb5vrYKbYGmuE3aK2BJ0xf1ZsofWno7et6FMcG
gxLqMzQfuMAOWDaqR7d2vU0xY85wdyCLeahoTQmTLgizFgMeGVBCM7nyMxiC+rhSqsEac5MN56xX
LIh3Myi5bBMYIvlwWig2aGf1MpwGkGl33Qo8ERJWgdWhLjYOP0jUdAr9w0s1wOuYt7M3FXq3tKOK
hrpall354qvLK4cvHuqr2vfP61LD47CoaA3S3uklG9GcidkuxJDLzhzFTcm74Ve37umJ8VA9zsXy
0IEdpRbk/FoDVuSSQyx2DmqoHbFmnTJNGG8YHtsR7dRyDiWUzxO2skoaY5oPB+7SPhnRr8NT4uev
weKGEIC7uho5k8Th1o2Ry8Ggi2h42bw5t1jLDaBhESn+z+Qs0zzzeK4m2AxdYy4A7zzNyyBpSJca
FaxlnT/YBl+ALGeH5gfO9GSEJBARVntCHEicUCntZOc7YOzE19ormNg7MEquNYvvxiEa3Fg1O7Uu
LKL7QMtxnk8lYLrm9NWphsTeVSJXfI1xe1jWLWIpFedVAsB+188hQIjW1xtTacPbsT1U3O2hltR8
i8r5VI8u0rp9cVIVJhRzfbac9t7fcmVvVjd+HaI6rsAKAqqqoYhe1kstZx9DXasOaBlm9BYJJr9m
89GsK1LYTyo7KeEekzLKjjQseIX3EDvQrhGeT2//gAkKoyOfoh2uuAut74YsiUsqK0p3LTTl3A/0
mNEo6ivGk4ftMV4WK9xrJpGjPjR87fzprdY9yu3dyByvYXtKHdMT/Ebwbl4ytNYcfsJwgU6S21Hd
2bVUjerwztXOabteK+0vTdnTU5+vuzOCSu9U9aLA0BXpBJ9f8MYWwr4rg20xRkfNZ0wigSdVNbee
JX9FhqIK/oYUWSAwjQLcN/qNIigvlJYB9LFQ0L7URZz+4Jek1BZHDnZDcA26b7FaQ9vc2Qtd/Dve
seF3Lun5D1uCU27liPI9daB6aY7gsahnKuWqrHipW0F1yP093nxMloBzRjcaoKBMCs7C/ZUccgs8
nx2ux1mB5i9PGDmCDGAIuAQmX42SSeGXB3XK70PIn5tiix04wgcxAIMk2JSdDS1d0CCATokPPyF3
Pl1Vsn0TG6zuEFijVdSkd47wbftNBRgZqdY6E3lVOHLyvv7eYPSdu2pbTrcWQ2myP9+Fj0b/Amgb
jawOjww2vKybLofDURwTKr4yejjxKoke5rYBaAdRswJz1O6G8tymWp/87DYfNT0/TPbcgb8G2cuw
AYBjZLAsRXDU469ACrk8ZyDW6hRA+J6O2NBCA0j7EqADBCW7f021Er5HAXQG8kMEDXKzffKD/944
F1/HhZckjLzXQYFmVhLP1XvFKaW4AiJYTo8ttYwQ5jR1Siqow5hV3x0MEia0VyNKtNUX/TChyJzC
aeyfh5eoTGCTtcqWflbJ7K3S6yG0Pj8BgjbRmZI4diZVyRda9lpAX8x1VFB6ibRIIAo7fNJAJI6p
6N6BoVowUF4ifEIW44mnF5zn31A59zAP8h0Zecg4ZjFsgjzWHJrFBPKPCmhTq6mzr0pLpYgB2VYC
E+IFSdcvuD5E50drAhoN7HUj/8N1kYAhoZ0xjIXWBra24C+wezGpbqm9V7fKzqcnLabfeUj+Menr
4bc280FTOe0n2VXQYjibs5os3RJVYGvzg8e0tVrIwTxyh2J0q8172fAOdes7vtW9ThzcTjypt9zl
IslbILdD3WuvwEYfX3S2oSdQXg8RqrIU0Vd+jxudlRxSJgjx0pBby6M8t0V/hJ+Mv7mWlwgGlR/n
o5TEa5XsOEcg3/sK/SjI18O0NUSSdpzCXVkxQ857pUVEUfyiKf/akxIz76qlH8jSFJjSE8ngo+PU
esS4+dGsRBInRd3v+1NyrzJ/TDoHkaidbjof+9k+G6xoosNoWnIGQ5L7Z9NSAkhBDkpSp/xAsXk5
GnotOgeeQkjQa300OmLNMNsU0RTCoEiaRSoJWHxOHYdo/stjuWuGN/ccJqWhmnKQrprennWiZZ5I
c/oep8qLjbtzsTbcEeS7374WG3J2Y6PrluHIhsfpDg9VuCYiJP5vCiZdLM1WRliMlL2PAHXXopFI
v+PY7KItMw0mA/1DFj+vwVZylMZzR3apgwc+FSLMDnM2/3fLkINNmILOZrV0bJFUx6xiUTJtmV6+
qR4lJvaBRyC0wqBmX3NK0t8b1JgW1bNx/Vkr0NmvqLoTJAvqzAbWlffZmGL7O+lPkCW5XfHisqBM
FypC3G3Ze5+oeE0O8E0OfLwf0yNJ32ffTF6Komzjxe4NakhBw2OLH3I45U/HGLGLO1kv+PBwQ1ft
O9DnA0nlntSQZhoymqovoLXyPQEkBUT7vwT/lpJfjELa80JDSbcHLYH1yjlnQQ82SBWYs8cuCXl9
Nbloy3bKk87t148BkwGDq8Co+zuOm9eSn/5WqhC9n4oK7VAQ4q2b9u0oPfj8/tckycSA71toaZmC
/SEMo9gBWpaEfcHn4H+tsSwlryfG6kmiky6FMcndUwLsFch6RmNXPgt0pY/QgWJQT2uiWj2yW6NR
83SQECcLvu7hCK/EL4nZejjDCB9r1H8Kbw8CTeTu5JkPGU9/FepKncfs17fBYDkVnS0G1akv4Y7K
uaINtQvxXfMv7bTitfrm+lw4p1ZFgRYu8vQCy5eRAFcSGJBDun1h8wsrCRZJEIOsbJ0EIdkeriK/
nraErZkC96uaOtL2a3HtH0k/mVY85631tPq4zSUmwIuyG+ENwVzvC+ist8uT87TjR5YdUCLoxhN5
F+/R5LLZFUQbaJKeJw8+FAEPQI9zOMwL8+7HE7en/oB6eADvP4+mU1l4e71pQugSKlislTKVAqcO
ezmTz6bKRgdFGWwjxSREP9CLEegLtYX7m8ExTaG9hmnJzFr/8u0if74sdrElBaxpKBOaBn4l91TL
g7J0Ps9keN8FMhWUWmra9eG3Qh8cZjCI+fv9MC3OPaXXX99TttX45MP4ITzqu3CzCJF5hhakiR1B
CFuwiehEerTD5DmJ0YH7tyt23ZlpHMD4d2miR9vMj977dZVvSi2V/Mr9jYbli8DERqdNKmK3Hg9L
mIshuo9xIPFIWjxVS7yktUP8+E3X4s+xask8gAvs6yOaotfkxT60VhQrr7jOMPrwQ1vXp+mqo3Lp
WiNkYYQkFbjPqBJuQh2fy0cULno9BTYLmte20E6FVHQfyR/HK/fPgUTDHCLLj5n7frgqkdtzQq9i
wtZQpsspqtybUzvv/m3TtyMJroTrI/H4No0BucCsQhhQ31P8i7HXTFgsB+Kft/5db7epP2LMy0YE
LiqCg1cK/s1FlIt5sRz3x+tw0uCaF9gt+CZHDeC+FOu1T5+akHe+OP8pBwIXHQBAXY05DtWzme+p
mHJAZkAnnJOimKayAJVRXi4+BWaX98vXH37qf1sMvOqOz9XJg+CxOvU+UDh/A4huLEArraMKW37f
5qdWq/uFjwhEbEa7ylQfB8Q8er3nYzdOMTg6F1EQ1AY4G93aQaTVDCl9aPs2zA/CrdiGFI9Na8zM
+tXeDHUf0LkAxWjasibZFOfzrou5sie9zI1QrakVuvhWjce4/VNIMOfVVy+9jec6vugo61qseLOL
IdOkwBRebDfDOZIzD48TQJNMHTnFLIlbMmEKPZ6xra9NN+RxTklO6O5dD91GSa/YkKhBHSnfSYHz
JZXNWAkmmJ90QB5leiH8knSU5qYZgdVh7n6TL7C8MUWqHO9ni1YKTNZ8Z/6nwvTSBhClA4Dnmgke
oA0urXNQ/InCR23p2AMIfPwNwhLzOth+GldN7onE+HxiQlPRobVnNZwJa15UKiq4giMaVGWcos/+
WHiPwbuNsOQ9o6f3ZSItASXhjMskCQ4MArX3JxrGgYd/Nd6XjUZESttrPMjgF0rMEohRJgWYI9sC
rwy5wEbLnInA/E5EWvXFNU12w5wP7lMncLNkyG0S2OQ2IZSLpJn4k8k5pqCRQMbv7tgbpmKj6osL
LqbdzqHNaQuLqZNT5GFrwIxAzbzaaCzyEjfyJCyGBMCEwDVr8eUYiq0eQMeT+kMI/9fe3h51NzYi
rse3pPbx5h0c9aDj1aqcUIG+CJD/1x56e2/vCts35Vhj3SAGpzgkkBV6Z6C4jJK0pOxbYWqr3efG
mLAyHftKO70yXXCKU4+ZenX7B9m2PimvD7LgBSSNAIQk/zNaH9VkyA9iGA1VJIlKxl30Zlr66OYP
F9f6IkcWNXnSVM5Nq0v43XK12Ir/VXUL6F/NbMbi2UdoHHJ5uPpn6PjaKYoxNfJ9dA7qNrAJM1uT
hqQHEetTpdwgn+kuDFGJLF9BgjRXe2cshLDpaDcICaotud3OAcYp3YtIp0MPb0c+M6MODm+H1tHD
XxZYuuU62vd7CFDh3/vJVg/4fEtDIME/DnNQI6THKpEqOyvbMyZ0+1PfDO4vxaTySXs2Vb8ALy2u
2yqxQmPO+gyD43r5W+wSdgT+9rk6nfnaCe6FcolPJI7pJFpoH5er0eHxR2TyQcOjF8faR1Y/rLRD
iuaKf9uVqd4miJl6BPZcX8hl9L/1PyUZheLUWOKCQPRQp6bY8mnHxj8QlwOCxGgsCvL8udU89ybj
WovfEU9zyu/UfzO0TFAzL62OThFNs+i9+hHkeb8H5W9GqJQWu6SowLpyOFD5H4SrdzigY7Z2Um+p
MMzkka/XiaTXsaY3lyIOZX+5924UD/7ZUGeof0S6qZzTvXcmEWfMSm7/M6PjV0wa7xpO8JhBzC9C
vlq7Ffgz7F9Nsxsm8uObFLbh7oGliNia1HdPXJOwpNuFLlEbTDjsAqcHzb3TWbEearUywbf4jFoK
nSjLNVET7G4WTFFkllt8uDOzo6Ks1IpUxGlTo7zcFGd2i5YXRtS8aZmRZMMCokc4zgc0/RmfNet7
MCxlHLQYItGmYGn1eZjJ36x2JwbFCAMa5gLqvK2gSNJaE/+LRQKXjl0ZIL4rjRKYKeVikmikR8Ye
WePDIXYSDRmkp7PG7HYehIVtF/dqAufEYa6PZOfYm67JOM+mKeHTtcsCG68FOCbclqpr7JK/W4Kr
cFVwvM7y/JtXUNX/H19O+NZlX6dapogTiTyjRU/8erEgXWmQ0mNQ0ce8azhiJwRUaAd+bhLRzhAg
+kjznjIc8PJQpaNLwZDb/IwDfUJqvvFk7o5KGfid4gjrg9Ym+sn6GHGoigTpYs3we/tZvJF2ZavY
9KiHrxsrpbKdVFVFbSyxE7DuqdpBK2Xhy3fffoMhyyJBOWVDQ/KbgZ34oByAIJdzFF0LGy41QNfo
Q2ilZbUP8s6RZyhp8EH5LPG7tiYyVlX/vJ62GxXhigWrUvlx/43kPyAGzc78NpkxW9Kj2I7adrvO
tOp8MLlYJAvcngYFucOjp2sX5SJHtr9CP5BcECDoStMAkBuPn0KMhYXfPh0oc2Ns0n4KgHRKCw2d
4+p0ByqcD3vf0d9hOL3iynLMO5RPXORqpq/1gGQMgqXxJn/B9R0v2cOnT4tfSpTL89tJvEEi2rd7
IlCSls/KKPxoVbzCJhhxTkaRzCzIycVCXOqf8sD+fBtGaEP2NRYuR9SQcpRydnFCL6eSIRBM7sJV
dK3fE0vGgAtRILrYITiNFB0FdEMKReioCUmbuPY3+Dgh9YKfgkJHJMNge6UotJp6AN04eozq3r4H
8MiQSKupprZw+5Fl6ffShtDkL22GAAv5j/h6WOh1sNcWj9nY1mdbHiDJYwrTPJjae03t36rBs/I1
FyWpxX7OnQ52R/8na0WffCiMqvATb608bbLzYk1wu1/36tr9ryMK7gEdQb+OxSwUAHKfjYtNTYg+
ZYcopaFCG7MBBcLXE5jPkK9JHGr/OuQ95XfMGPHaQuPiKW9HgCzV0NXJ/i/NT9t5wAfME2I/qtDx
MVcetB4vKy7Vp16haLxNridlDDI/4J2ldQ3Jf2yi9d3J6msxhA24nHstpoOllepEsktVZQN/De8k
b0THFBd7sv/HqseBkUnUal2gjZORu8EaLwyeDzxKYkMGKojMoIGo/ad/gd96jN3ssUzVbJNXDVbC
oYp1kS5OZkKe+eua71aCGqfDBvandiTl2ZJfAr7pVsncihutTS+mwCj6nX4H8YSF5/Dhe8FHSuxT
kk8ljtquXJ4KKoPwVciC70nIEkEgdrjjjz07FmC3Li2E+9H09fiHHNoAvW8VUUsJgPUg7ub81Q6S
80Qy1iCYuZ+XDcFSAQeFdlDUxJc6aw/o13hakW4RDd7zVQqebY4Ldkc6kuYa6DVxdyj3xBeeIABf
+ECAe/6dlUHdNjaPZf/DyFdl8tPDxk/Vv/2o5nu0lQ9VBF/3Y7ZAfT+evaoikt2/NmhyRfJznKC6
KEqbaNNuFKJKXGpX1BqIV4yOT0b3NyOotEe1k3D/K8cTj4zPfKmO8V5+vU+KXrrsHR607GFZR1F4
pz7rEexIlf6pmdoA3ko9iU6szSF5YsfRuY44YTEMo06yS7oElht+4LuTkzoSg85e/fbd0L3x084U
eQyMZNv1rcR4VophLEoIN0jqMay6SiP2svawLuL/J8vYNxHOwhRitVPoED23j8kNGRDVuWml4QPU
sWZMCaXJGaTvciD6SPjGkACvrFB32dctLaqroFuXGoeXIDmmFy3eLSf+mNv0uUUoNO48dS5lK2tP
HjF6nHHb9nTGe4yl0O1pL+GyCkGfBCleMzwzcWc4Z0Zu6Xquq7xg+Y+6VYxGDTiQpVkBH+FNOBKN
tnO0S3eyzzGDV3myS5UICjcjlNYyOgRGvpfbq8uxt1g3dGcnxyn3+TJzjYVxmbYrh5jl/w+EfypC
2ch3nwm58UiPfPa3rTaetR01tAIdHgp3WHFrX0QFWbsQ8SkhmGk9YRtETcNxT6r016D7H7wHz1r1
ju8wyUujEAaLqFhElZOUkTWo5IKjLpmaMnrEGurWGdmT6p1gh5QQMopJh+CU1BP5f8LSNOPUAXs5
pK+LRerqZxgfxK8Ib2czSp2e653Kxtm7Rxk4qp23PQzzrCkTpqRfTPJcFZWEQXvqnFchFxzq+68J
ATFC4EkfGSrCLtX7MCFpLlndmSBqJeTW7LNRtea7eE/eKomsRBTpdM021ofT87OY3X0vVEl5t+mf
BZaWpFsUVJK3TJbBByMNh57OLQHH7Vycuid6ClWTzEHxe4+GPe47JYajmTxhY6ARVveqQl+4mwPw
Q+3fhd1mUbD+OdcBcof2ogYYBt5vNMteK2Oznexx/AlBNm7OYfLDnXU3ft3CuJMOumXjEsF3Pc9I
oL0EKKyy85Z7ebeVVW5Rz8XRFML+DivVK40OvwHQylHQCsHYEzgvt2JRU2a80vqANwB3OSGDb8Tx
ojq2uGpfN3b9Ri8oKxN1xvhkBRFmGsuTTSMYupWXW5+50Btgt5xiXDhnbtzQa5o9wVJGmSeHQdUc
lL333icX7q5vfCYYmCdZZMV4rPcqpk1oU6yUEFUyFmOWHfRT8xgSW4Mke0ptp3DRkkPC4ssln1mz
2ibsfqeZCqzkPzZ4QKr8x6H5PctZxa8eS1/ym7+d2yrl+0U78rjjXvvTaUFDVMaY1nlds6j4FzF2
Ik1UL3qstkyR2ftLkZ2vow3+AYvrhVfGop8F/SKeTLkslbJzC9PnBX30SDAkP9K35Gm/8Y0WJBOu
IhwLl9AL/H4xRr8+nFItbxqy9cumaLhFFa5m9DxrUe7EVQYHpsNa8Udyg68G/Sv5gkgb3xb7GROs
XfX99ceyCJgGwHv0GOMZ2B5uaM/iQFhRsqDcLkeUic2bsNaKPQc2YMbROHASdjUBwKiJWWB/xfVR
1zEQJRoySdrcDuloILugGzk5gooK+a3RiByDXOEluzkG5OjFF8e6dhwXB/wcS955WIN2A16wkNhv
Tb3GJaSXA8gdML0deU4EO3USJU9NKIGCK23xE/2FDtteAfT4tXfhFk5MwsfZS1cV18eFVfkUi/J4
CL4gumw7CcZe1FFj6t4srUd9FJBIdavU14es8UvvAyf5k2W4ouH751bqbKkBFSMhgO5YgoD0u03M
ANu95kohLrCRuwmmRp7ccBt8f/UzUTAsm4ZgMprlF6Q1nSiAQi1exaLJboq3JTaALmO0mduMiNzz
HmpjYxRkHkUItXPaWNhOppunq0MaU5F1/MrLv76c867/A+azyFdRi1axwpiN+PfRaRH2Oj3kpfrO
ry0JC1EGPaGiyo2CTKOXG5H6nrgTFII6/KU6guJ4NHabX3f0h601nqhdDpo3wQo5pch9msF/Qb3y
apb23QdNG0iegpI04abb+Qnkq/x+CobVFdlrQjdvddOocGwo71mJKoesdfhx9SDGlAT6uM8VtGIo
iEYsJW4Lfdv+Sz9XOWL0HCU05q+LcLCZdlsOn111AD95WueoMB9Hfsi/fD7aPJ1T651J7TOG7mAH
Ic4kJoMgcqRNe63hgJxDgSppN1EqCLxpAPFLzpqEodixv9tPiN15sqEnceJRHrY7H5ah8ZzS9xwt
tiVHtOR13Ezqb8JY1hEEPSvTc9PHh7Xq/1lW1KG0hhoZ9YYCeb7NbCSXmJLD67byN1g6658VLNY8
bTKExraBj++mVaAcxd/M7H37q3VLV0js115eEQvX6+yPIZ+QHk2vskijX3JhWO6JXIheSTBzZcG7
yeEzxvxVCWo4ReDyOnn61D2SASnwEhpozCcvf/U9FucOJYkKtb6oz7lhSx8BCOA5RSZpaAdRI14k
QJfII6fuFAJf9LEwky75Ecnuw79zAmJ4RC2NwDIMpFIOzSdTw0AZ5S8P8SL4qykwK5m8gBcRjQLi
vxzh7wkJ7IK7O9qKt9DAWD+rEIjgkTO3aUbTGpBmSZlcRrEcS39Pm7c9nx/Mpqastfs6vsUAHsxZ
xxNIj/zYQm68gOwbcFgJJxdPUNjB5T1BjxaUv13XM+uGsUFz7ox9B0o12dlOCfXsPtBN6+nzs2dt
t34+ZK6sayGwKYeKzfiSBT6GcNSG7nDueEMg2/aaJAv2164cEkCwJECxcogo/MhcHhjo8pD3ZY5N
th/b8v4zGUssJRZfaAnXXz9AeSAXSpMQgDZEltwFfsms2HgmCuZZyaJUp1s82q2KNNqLYO2PTfxR
4IMcOsLkqZDy99eOOkb/rPSMnTPJtJNS8b+xGEnvOIMvZl++oSEd5sKQqLpfna1ny3/4n++/qL5x
nI+QfNDLXGndFuDbiB8+8hq2Ez8K/pxkMgD62f4rjc/OxDIKQ1qxymyPTSaTtVq6a+F8/zstmiCF
YYWsaFDE9EPjFVAjvDLDs3YN2CyKXEwuxPo/L7Dn+EDjztw+oYC9PLuxkNBA2dnNzupWRFxZCpkg
HLahkrOB/gy5hwrT8zXR0CeeG8JFgQFiZzWRMrvi8S7wIRRcElehQi8Jsf6bJzohM9VeX+kTAS2F
o9SFowTPeLSTuyTvOAK63jxRsL3d3dKp6wdWR26LScxq6d66VrYeThAkiwHHRPz51gNs7FLs/gvO
FZLP0A7r+CEXMO744WYZj9jtqCHn/yOlM7gP3sBom5J5vO4aJlC/Qy2wYDxBKeRKD3b2gcnNXHLz
McaBk2yRpawTxk/D/K1GsOap8hznXdDeq9RoNiNmNZBJE9BabgAfktCRVxG6EBM4vNzn2ZVB6Kjk
A1eIBVagaHpRt0T1ToXtJHtQ8PCklDHV6f0EnhrQy57RY0b70SFBi2c1m1684emzXpN/Zv6qqjAa
GUsSpWC2v0k+fnrQkdC2jsuk2N2e7UbXRZfP+tQbFy1K8Zy4qOuk52hQiWxkAJf63eQh7ehKVBeV
534FBWYeu6a4L/KItnk6NKFQQs/Vh/H0av/miDOme2Qw2MnpuPogXu1gz9WHefcf78k2VZAKU+WY
12hWGLXNGCx+21Yu/mtM1nEwB7mQT0hcme1bSi3N5VZtdzGYLCuOsDiRNDlYHmsihYGAiNfp3VYu
E+ZEIaXkYUyhyFrN1FKkOWv3GbN39vDCxRUdwTOQ93hY0BzfycZuStgLEpkCPehEX8/onnYP5bVv
O7928gI9/h/FpTblPm88ssQJqDqDbhRmLXoWKAYJwyyjICQfkQWEJthS8c74mScZgLler5GXw88y
50emapzO+U7EYYgGbOVQWKoqd4aJQFu1PMT9qm8rdQ/rb9dmo6t+rA5MoGKOjDp+W/K9Nemi+i1P
+IzlTDjeka9t9cJKFBMmNozuZSOWgKEOHrBSu5SJ3ZqLD7r2ihdKXlL4L+hCAYfoTzIvtD3b5InQ
ZZbbLf8xVXZK9GIg6MuYS7BnDSg4ZEpWzyNN8rK1jDDRWlqaYImO+87YTjpUO2Tlmn7vE4iELTVm
qGtLlFkG4/ctY4hpJM9qqxWIgyz77lzF6Qw4i/5OLOlrLikbSrbHFOe2zfbDiy+E5cffkbQ6QvpR
6Tt/HvPMudgWqYf1iF5ztsDrP3HCCqSkICsAfBVUZwaMflkSJKLEWx253QRo6n4uYP2yG3/n8MG3
FyjHaBKISW3T7rhZikTZuOMKbnFG4wqCYY9zDk2kDBhXhANg4tiw29ekMKP+ls6Gpayb0BIGA7pZ
+DjMrrA2+hE6QqSfzxIsoPPmS6oaWnM7GpdFXWaPvBZVFfNbI08U6xLkXFlJ2U5NVaQOc/kNyFCn
Wuw7FQbIvGMdWsemdNVEKqasE/yy9CIZ9J+lz26UQ2Wlw/ahn20ZasOewkGsAFNXTv7z65M2klK8
piHaTYILzGr9WHJ/iODhmC0O3yx7HPY7nTE1ZgqKHgV2H9yTgVIJyEVMFc1+IP3i8SKuqrsP08Hn
HfeteLyNVZT1iMLV9YtWa8VBmLZDwzKK5K9xsxGICmXF+Ojrk12lwF3GRbOzSnXuO/wfPNPdE3Qv
FTeefA2nVf1KsDz5nnwcgUEDq0Fp61WjRt37Bi3OFe66Tekv/fw1XVvUIZTInRICm4GLmUiIGhPT
Spe4vXz6E5x9A/8DHKybvtKiREjELi2xv27YoyTcOjjBiW0FfhVrkoLR4I+fLxVz0RwH08fMqs4c
i34fq/g8K8qqzq5jHhfoYaHDTiUbVOMVG4zmwCTcQhcJCviUsTN7b0l7ujWpCuS6kXp1OH4fy0kG
QU0UX00y8g+/7C3VY4N/CaMZb2JomAC87o32AB1jbCVZc/0mK9A9kQTNURDvoAaEk2MpcdAgrmFy
p+SR/EqA8cEXb+yolsJcWn+AoiaJ8lEFVdt+gEOuqSk7xAccHjfN80a1LUHlTrobi4JJZzmvmf9a
/fS8HuWIXNSnoR+RuEHcsUSKWa1vEr+oJj79/tKf86lpaAElZYvE4Xz0GvW+VaLhm2eGOtqNI4VB
/auNauqlDbOgv6XwBj80T+G4ya/T9nJoNP4owewshWFNAuwN/EGA8Y9NMVrlaFHLSGpcpk1gACvq
/2PiboCHciIg5ufokKaXMQxv72h7dT3+GpmLbi0D9NNuhS9J3hIwOx0QFrj+7/htI013fIDOO9Wm
bwJqIoOQevM4sSGhhEjk1E1KfzhCQqMU7Nh2MKglrmRYhU1KOkbVTuDx1ELnbWNuqwIfZ36+/8YK
ESnm6fRaK9V3dIsplAlPqCIU33vryPG+cYJ8Cdn4l5A8zBOZkT482jHt6uIAUlu5egzIOAtNQn+A
ScgG6QKPYXiP+CxirHBxl2oZhIYTBewmE/ApEHLJfKLBbPEWQ9VhMLlyr0CNi0kphsf+05sSypip
trFCj8UxCRvrcvqov9wl/CiSoIQZCrKeJ0XNXy/SEzJj7JJh05ZH3H79bnsQ4o2bvLno5Auvc8G8
iaGAfEbHZnSFsKXQC3+ACVRIG8hECIWKsq/4G5A2f3qIhsNRALOdFFZxGsCNaY6qRUxwtaUQX/AS
o5Vur2yAiwnWsyLz4UTQKZI3eqd67YpsexP6nLYhY9HO/04bwD2CdzzNIkexHOv0KEqKfkiJ0vE4
dIN0qshcR8Udkk06/fANY8e7VvTQdyVaPqXAd5inZmVtQc7ddCOThhapVAAu4csM/P3WZcFh1u2B
RtaVYf4YrusrXob/3ToCDYWeD9FRzJ60tFZtZcuCpIrDbKhIbPG78v0kRio1n85c76wc+qZM+A3v
/SXVfsbVdfSE+hBIsimajrOLcjhY9YexbOWUq5LXrWPu9yK3KIIoINAatCOVKTkGnGO4ZVw8gPN0
1HpEYtWXFpo5hDeytF00Ryj7CCom+pfTRIIm9uCC/zHPIBKu0KnwrtoIo6qfhqW0IBKy13AbyqAg
QgD2lYye2qdyDSrODzU9hRdegUmdInJ8C+j1LJ8mbRx247c4D8L1i9G6g4gHrhqE2PhhvHOkERpU
T2HYbj17wo2RTBAP/3DTZtwDF6v2xgwXRdfNRXVjvdzeqHr1nKHIffb3gR8KyW8b+HY/FG1BfS+i
mo3psAHNoTBU7p1muoE+MbDrtlExnRm4Nx0G5kVJ9vSKwtCC259bLYQBIRGoJFfSdwxQdycA4ZA7
saMdbGiJMEDleh8xiATyD7t+9A6Ng/vItPUkHgz3FMi52P0NZgYda/UF0X3HnZ4+DaY3YSLpyJCT
EGsHmQD9e82zG8IokdkflroPQWh7P5u9fmzllRbWsZDBmHSYtb4bRvufWV5lXKVgdVVj9NkW+4VO
X5kA0Yb7Zbz3Ib942zJL6yLFHc/6l9R00sjOGSSFQgvwBdwv0KT9+rIUVAYY1CYZQ81tas6P96Oq
mqInWIXdW+V6aJz/WkVzkRpm1g0TC4a2fSuqRyXR/ZhV4OAF/uClhR1Y78fgtfpUYPKDNv5rxKJI
2+TmWLA5Q5oviC56BIRcc9W16AZKzpNG+dKgWlh6UnyPICHhtkr3gdNh9+YwIfpNchuAQSViemAa
1WKgQsI41x/5tFdR/BAVXckWEzKmVpmpvALbGk2nFkv63V0GMZGWvB4cmmU+ureB8f2gQxfh53PM
bqi6WwKhjZCwRiIB1/If0jHPMjA4wZgPl1Ur0b98+jf+32+U0GCmJ70t/jhV3oF2iEC+IFuztRcs
u6Lg9nwgRqmI2DFk+Oke7z4cbKCdjgsIQgmkd35Jr/E+AqZz7DP8RSxSyrxF25tx0Y+BxA6s9C3Q
mO4WYu407uTexRcvzdFYdM2ytkCavltQBX9hQ7l4u9sSb/ZMaI9DUcdmIICe8ceUihFflp8xcjKd
JGkK/j0iMOMP1YGRRkeZPBTusj19HGCyx0JINgmPbqs3KzrAKpeN4gzZWX4kUw4yvq+lr5Kzlf2z
QGVxcU6OoTMKQ+H4mlc9QR7UrXWzEY3enzWvxYwtUMzp1E9xUH1AYyCGDsjbEh5g6kXUJDJsCD2y
u3h/Psw0x01RGnchXER6z/zt3UaymRpqKVR/0KwupuQfQN4Rno+zhqdFHwj85tqKTat1HHHlaCxa
MySmC/UHKmWCiBYycL0/HMfoQbSBAThiQuDbhinziakQ4kyinq7F14+3BAroGTrUv0hGPs0nb/xp
Px/G5nUFgaqLo1ER3fsxfLWX3KhFYxQlph5DRM+vaBTglKm1KJbYbnIuB1nrF5X8GjUNVm/lCpYc
HWqkOFvFMVRuyVon2sTSR+a9SFh5UOt16ArMPqExq8BXSk07EMqUJsCbbfy+RF/q9ssOxh0lreW3
jiGMex79aszpE772eQN2ND9MUan11oqXFKgmDaWtWehZiAkNw16xOKRSkN7HOAhmbLXwNFvSwPyC
0DdPtfm+gETtS24mfbaLXykd7BB2AHSU+ar0wKZmqY8ijNWTfs4XaBqMQp+2wWp+l+tYTndDXwIE
F9k/BU2OLExz8FvJ3IJO2Akos4JjbysMlMs89NlrsmfKb6+UctqRF9V44WtGfm3q4IPMRRj6E0TQ
seKsMoQlAbskIk9eD55lDEKzO6io8dnRJqSN2dQtas2NBGHnzzrkpr61mDlJyeDZROhHvLaQHm5g
NLxMPnVIK+vutfhfvqbwbFs/98ck9Puk/eho41Cg5fN/V+UdZtOZCLEmjHKYX1QFIavuWdnhBZWe
H0IuKxLxNtK/yrTcOEYF8OkxXDIcyaKjtia3nj/s96KPEctnO9B7ZSUhFNZKSwa0ozvN3XHjDd4o
lr2cvke31tS1yb829tH7dN9GLZ4UQlctcVXaTaisK8CAOy+KiKuAQ3zVqpe63BN70uJlslEKb7ol
LqM7gKcXjq+fz7wCzjuWPurpER9qxhirzFwYUzZV4QO6ncDTWv/Nh9SEWhPFUh3PmADwU2Dz0XU+
fI26RRg0wHwiurUlg/l0cq1+U10G22dq9EBWi2wqkKQXXr7wlMVhhs8koQzu/OSNMfEUDSuh9hfR
HBJE1wzKvo8dCPk7EAlHH3xg4fZa4axUpY00ej6Es9L0So6HE77fPSWtb3YsLDcTUP8P72HiiyO2
84ElOTh1+7rEocvQtS9zImgoJ6Nf0PJOaoErQDG6NL39VIKf3+m2Kv2nkVhj4vnsDah2GF7z++WB
brrGiysI291de+TU//aWOgkQk4eBeennwhwKXWMsIxPrnyWasG9pSukYgPqQfh6aaerQVe4xowVa
+omIa0rGRkNnaY940j2E6UYd+IyR9Gvd1jbsjQ/iOkqlU2d6f1NTTYrM2TAtRH00dKw9PWRImT/L
FxZJTUSYIBVEdUiYnMzxEYSckmAY3j7Qeos3KYXwYtbdjV+6YOcLxUna5eAOxyGA3tbyT8oXywRU
Q/koZFBOCLD/UYrxuk8IiyrwnOXqDfrxLo7AGE+V9aVvGxP2G8hCrHAgMbMYbcRGYAGQ7WPbzuiN
F7M5wFf4zB6PJzpYoU4oZI4+m1ZK9MVIpz9pc03cdxSFliZj3HXR7CUQlP6Tb0pPOTO/Y/Vfmy3h
j2+4IBqJ6oHqN3l5kVlxfLMpFg+kga3pJVMxHZwAVquQgpa4837NAPUPp/TglvAhHI/S0fvYqpgJ
vLnDivVs6m7tw3nNS0HKSId/atYxSsvvtdTW/9oNRkv6UlhvHDKRXU7/KJs9MSi/oeNDgZk1zXHD
qWk9E12O4qSsjPTzzobYeoMAoBTdCzax+kKOw+9f9Tl4kl11dPCHv4A0i8dhWFP/P4sbK8+EojNU
uqyJMPe/jnhs32kc3RqoLmdXd7Q+AH30zLUA0+PIkTNMwuSTA1wwCB7hwnLDFyMiKmEgrDV/FwUj
kAxQnheNQAAKbQfqgc4kzZV2sQIL/qF9GIKC88YKkjOzjJL+UMcWdSgGC6qGrP7gq4dXSTULTgWY
DlKXdjxp9/FiguencvqmQhSolUnogrr3I4zMbGntNGsc3E1qFYCO5vQ0N6ybmMrtRXSZIWppfbv4
OVgnPK95u+AYitRCETrwIWSGSM4oyNivJSgtYHi7ODWtu6udD+XSTZCkZfov4YcVoGhgGUl/nnLo
o3dCx1aT784x2cZLUBVTz7vCuvrbGyd2Gbo99rHPO65eFendZoHDWBWwgHU/5w43tfeL7AnffPnj
3MLfAiZnabK2Qk9RCqQ892nvN9B94M3BoKAtDMDXH4YUNl2RzvxewDiYu9Pjod1uhZTdd9TyOQ87
kzGacJ+HjW18uCAsHHKunR9ZB5Zv8GnA6ISGJ7ksfB+44y3oumlT7GcsR4JGlPLYX6gLTJngB5CB
ZVarARaA8E83W7M2LZ1p6iKnkwSkaD1IYyMgu2vMwqiSYn6K5trimFcP7gZlb34TAggGX6xV5w1d
9D7sdgUAqax48KH99kcRHvPaGh9AXdiGFqSfQtt4fO3EFIoyq/bZUe7vCdT/8+UZBWvKWr+e6HX6
0gnmMXgEJ5v7Ypp0PYDmRk7PqG4idII/wl+vfJc5Lg1VI35LkGysOmCVtTtN6zbkYSpZSSGJs6ns
XlgqltVGf5U/q4HVar0fLPHhAkapN4hRDbw6bCK53azmE70Ku67kdAEkhq1yqj6/vLLm/YfLBLLX
5/nGaaEc8U0cRuNUUYhyzXe0z/mnPIoSGjk1RWHHZA/U5BF9xVkJO3JpuwsMERfuDphFo0B55OTL
3ktm5Z6+ky9CAzBOWzEQC466EwX9saDX+Sm4g0tjiSUzgmwr6CFYJZTuYgSj6drahS7FOukd30lj
siAQDKqlctF1N2vLZpELrT0ALDd8Jy5Kh/1Lon2cp7dEA/QmrMZvA2v+7QYeOYJzn3i63LFsfaXV
vb8TaA5TPUDy8GjErp10Fnj2eC8D4CZeitEOPsLi3cTJInG8QGAtHONL11R8A13Pig6a4z9PvWFS
rIrrcHzyKl1zv/J4X1S6CqtjMnddBpVRQ3BHfZgROyVX+wmVEfHAjUj8jzMSv2cvzH4sMYAZUAHi
QRIFZIcHg8+6RdGJnhKEcGrZMxEcP1SuP0v1KqbTYoB7HAjHTNr99CADStHEEDyq0LSSraBvrPDs
7CR0KH2W1tnTx630jWkIUx+Vhz/SwA9yBb1AzKT20IiTaFx33VL+8tsaU2wpBeooQB4RO15sIBNR
sfUm5Q5UAAvOMWEDGCjutjJWrhvCi/rEv9FsFZOf55RXVdJlynhOyJgWCwkH2Nl3BI3Km0+kSVd3
Ckvad9n3vZXW89fwiGZvlAw7XMALNLcpbbUP4t7v6+SU2l0ZuAIrP3EekzyHEdUliZCn9gXNIxZR
dewjzibTGNd7JiuoVQgdM9I8DBFbhD2UAczJutvLPQYRW06dTEfZVd6cnxr41qUoJj8dE/JizLZB
pKOaTjfXIOHgZaOQcH7wUxle0Yp8WLTgYjc0w6DUUyXOxu9gg/yNBnsKwhBhimRP+V/0Xd6CIcHg
pChbptb/Dm7AL1dFJkSo/Ud8wROABWCTYySyS69QFTbeq6LUc9CG2HQhVkTRviRsVeaQXckHV07s
Pf16CmI7XRjv5iGcz3Jjjgxp/4qTKDf74EYe/Y+LnNXk5OyVzXp43HrzfIPvwKD8jdGq+MwUL3Wz
DKCG4wDhAbV45J2Hk8kRDRSa7Bo6+np33fOqvPh1hC8F/WWlsIjCSn4dZ3yIW8sIDMpoBFx24+u9
GV4L6f04agY6e70Xcj9yoMP+B3mw44Qvp3Vwn2Ze5j7B2ss1srr7X3PmzU4lICO9Z7rXNwWhX/5A
GE8aAukVR88KgEGudEP23hpVy66U61azcAu7pJaAwzBh7GZEVgNmzogEFUUY2a1+PesqnPouANmS
7Erl0QBcbjNyVLoLclrH3ruJJ/QP+yN0vZEU/1OKGih3heMJhpJzWZVn9d+MSJBsG5GtmjXlHyNM
bvj+QWWEPA2Gn4zXlTzwUchHIB2ICd6PJ88QLwYgvnL0vjO0yNZap6/PUHv4EU1PAe5q6k8ZAydU
bsGdVTAnN+uhs2XAAGH0AVN3U+Y/tE708wYPXAG5lgyHGCFoGo7Ko1DLWoBMYpCY56NtEhXuIqMn
oHoPkeaBmo1wb57xC62I4MVC4W0jKC2Bh1iP3oGXgBlDOQJ29GHHvc/NMB6FQkTEzRQhK5xPkUpH
XXjKzq1kYc8ugxfEe+GKtbepFc0JN4FPObrqaewmv6ZOl9yQfmBCChQquhWNVho505xvjFw+fLJ4
5JOeF/oeRK1VYxylFA0sJ4DHh9+VLjSVWLOG1jAbNAfSrmH2Q8KWBdQklU+LAziHWPs7AxAv6sf4
J/kyPxOplMa0QPPDfnhKC0bvm8y9u6/pIO6GoL2VPX7F0fY3o5ZUFl2MEdUVr+n2cWMB2SFm+NHB
RPEuD51ChfWp3+q8MfNubr5sKTl29v7Zi/MmfxVhNi6h3MS5eM3y+mNVzQaU5s8YM/doRDfHxACG
8fBOt50DvxstaGT3Bx00x1rIikdt8Mgz/et0/YWzlaJJ9ibeZYhDM3hlyxLfrAMMkiB5gjmv2nFe
xmjaFmCxc5LZ3AJR9HXJbnjV45EI7hKY5Pdx6MQ8ccUz8RXnXTF9/+NA/g2jmKqHbVNBePoDMNot
whMolgI7Os2tgl/UfTl0cJMEVOivS8Z4nV6gRLhd1nH41zVNKo7dMpIF+oUVqcaTdATweGQpuubg
JziFp5UUtYDhpBMnJvj/pPnMBZCJ5Gqww57RV32OwOZSIOFbqovuthfD1Wq8aN0IflkGM61U5EFK
a061xzXzTx0zfu9AI226hLUCvE+xCCYYjA3kvt8G2pSS2xAXdk1a2z/GdwwTl2a2nFreBw11sjDk
xhBDRbUyB8LB+TKQ07CtCGoPrudiFL2DMm54MmWveXs55qnXS+CrgklpS+Y7D9rdihTbx6b5bPbf
6jIM3yasbHiJk5B1zbLvxWgujVH7eHe3TBOFlk+0l5PFS/JuWmTLKp8/enoFsmEpMmSjOnv2XGtR
1qhHF6J/VBjgPVE7y6SQq7tW183P0GvdWaOHw1y2B1F9wV5faETAGDZKT93eVaIUtytfEqtIZdhI
HN0Fp0fGuK2/UhyO8oRCKM+DtrqjEYlhfRF9Nzgsl/0BVhMpYpzOJRKHJq386yj2qUpgv/yTl4pf
DoCqQ2pVUUxnnE3witseLzSL5BRRnzucLA2H2AjVAn/aqAOBfC5kOm+nD3mbqG+iQG47XlZg/GBx
IQFz9JnPGA70cRhg1pMcKRePMCYnNqoTBJu29BOh2gPgpsbhftHimKDhN1xn0Eq8QS1Wo2/cAgZq
4gZxHSaG/tqpGzYiI/IV1DSPyiVcwN9saEEL8ySlqWHzt/z0ybvSJRBfb1suCES80jzEMnQuH3DL
nNlc8ZKwPvbi8JWtICAlo/SskNE/QHY4U9uKH4DduAMAc51jgOLj/wBwYAjRCaPtkIEqVna45IJR
3YcvfbJPtA/LEsg5qSbFKq0tQA7XVbwOh3UKsUG9PnDt8qpaVRNxwSuu25Lc0Moj4b8N16sjz/kg
qQOFc5bdCM+s8Zasr6Sdt3+NUYxstDVC+9eZ1Rh5z/eUmkiWrGwQLXVnvV+wVTYNx44R9rRRao6I
MBYnF4OKxtd7WgeoWrNuPpU+CfT6xZZRaDSiVs4IJwpJ5rtjeao2FaWFhA/ftl6S2qUk9hX9bHKu
IDXH/JrGBcuhgYpHKExzU1OqyfkfMVdxzJyiZAPPryhbiEopaqaKeQoGw2Wpwxw1VNj/KDYI97wN
q6D6+8TQaGcnfJlPMrZz2N7SY5jh/D+rrvKMTG/NZqOuUhyApy8lpEceLx8+KidMW4E8ddN1xBDt
5YgmE0D9gr7tgoU/AKVL+gn2H78n6jg4EpJNLLNyv/9eVqu8SAzdxLFQu2hl1hmYbwlDOxuNK+ae
qbmSoB+shCwq/eOs1NxbA9kxoflpqoDqL6BCu6x0ywLB0DuqBgJJaviH8AMQhh3jptdv+kMUef75
maBcLM/4YsLCDQb/fIsy20brRu6Vzv2jnj377LpSgCzv3Tim7TvwsTA9pSk/+aa+JE5OXMzNLe0/
2qaRLXoPXynANRHFcwpYp6UPIXoHiieIK7otRH7MNLV8OPiMBGEPbmAtIf2JHdhM4Go6FeIKWl/j
X8epICNs2nv7j5wvnK7w9RnCVZ2sEx0+r5NOp7wzgEHe5p1VDKIxT1EiH8YiuCt+U8hnkY40zf0i
Z0zLS2pXOLlEdnu8eFgcZ/F5xybnM6MKsxUkVtF9Uw0cuPCxxqeGwP1rBmNjH+YMGANsI7SWy757
pGGdM2UdZSZEPwF2m0BMNcJqLPPgoh8IzDTPysWehk8KpxPiZK/RpGB9LNFgYXue4u/u/qLnDNnC
vPwdWN+HEVydswtXO3VzwgqemUugHZyF/l4rkFdt6iZVClKM8XhOO3BqEeBm7Dwc9Vzxc1zS4L3W
KobtJvgTFRGhbZJa4sE2o7UBu5Rfrr51T1S3BMPJu7eCBYfwq9p3QHh1fA1x8lm/Mb9C+2BgraRV
8S6Vnrv8ofD4ELNCjHJhlsAwT4CmTL6eoZxa7mNq4eIpNNBLALIXlsU1/77T+9WnZqHFMbuE5uc3
/u+Jc6Acwd4C5Z5QJuuY/BKrfBEZ/jAdvecbSoxtEttPXhFKrmY/UhyfA2NkIjEZpJmI8RIf2gKB
fWOkWCxBxMrL0iWBBFEfek4iQfFI0a2nSXawq6xRghiglHoVulxWOb2Z6NsGWLyjFDxhuijIiCv+
mnP/pQ+hoZI8CcHzOK11oYMD7lc++Dex9hwaFiD8NslJea2kE32pG5tE8Av43lifJW/SEyJBIZKN
b0DhfRV4tFlIwPlCEo3NKHX5Pu7rlSrRxRI2HLfMOvY0lbwzq7rm6yLXYPb3RJc9SxT2Mpd/tpYE
2qi9uLYk23ouN908jHgAIlAgutK9A3IzIXc+vlx/JC7I25PAbmIYLLjk5sP5kJHY5HNYsyPF4lwx
1fc5hSF5RcXDGTCh5baIt8rvt09fonTpU3w38j8TvfHWqon9CKm2gj1zHkxoHj9jN3CYqITH8QDN
Ro5cEjvTujG3bKJ+iVxJTndbVCao1R1BmzRAZH2wbBFpsDx2ebtYkAqcKIltHth/ROyRonYjuZ7b
+cC9r3995n3KEQ/L1N4CEIs87iYQ9ImmQ5r7+PTFAB/6wBrJrRbz1Xl5HNHzuuVlCz+6E1bQfXE3
6MG7bVrCCStL2eUX2OuFQkzNiKvNk77Do2rITp13/CMpphJWmMfZ627ZunagMRoSl+pLhkbt/bfq
NPxkdlrW0n11MprSfMAqr1Bp7o5JRfwhcDPtgCp1f6OgEUaJ7pHqxxGqEhtuR1PAuFos6EvNnh8q
3UalEcD5ZyFHpFOG7WnUdeyXM8m4CCxRRJp7+84D9DjL/vEprO7yWBpsXyv/tvgYRrFYOwrbAYPc
ci7+lU6mhvmKXsQA37nrm9JyzP+PS27hINUYzhc82dE6izrFtUgrdAsiXW9S3clsCzfiKnrJ0Tx8
gXEM3/0sF0bRehOUBAxoxISxUf8RlPZHaPjShlh9aMjlOjZnCKDRseAxtdI0lEbxE/SJa2Vdl9zm
Q1TAh7jave8UDXZ5k3NVcAFZ+787BPU/dxlU+95SGkINUgFfZQgEIpWbRw+yu13JS1bIZeUsBiX/
WZUTros2k+COFoh7+jpjdFssFNkJhVQDxDCI70XWy46jbKwd5foBzFZ/HCaE6WFrlLj3nUPcD0vi
J3ng1Tc+Znsbq9jKwKXH0tHx5Zj0OGQR6RB6AyhUCma9zBZ1iSqC/yRAPFynPOZJs0Mr8HG04czX
ZAaM6nVgIpPlDZNsKxCNUMMBbCI7htOa2N/q8NYoTfo/56/KMgvmjdIKhJqLGgOQtxOh2Fpftkwn
xhyYZLPSb1TLVu9D430/HaJ2MpXGAgkB9Rp/uFodqzNuI5GwVtJKV3KCBRFAWHmCDyzzeQ2fomtx
j9Qk36ZvUuj2vTNeIbQMAMLvnx4U0dm1+wNKgkuI+YBg9aFoMtrVLz4DQyou3cNsfuefxPFbGfDL
2eXqh8PTy5vu5EbeRresJo2/JhKsj0XLL7UXGeh3HtLStZ4kNGBSwMcbeT06GqlEQwYY0e42oCG3
eZhKnoQG/vlQp2+Ja2c4fsvrtU2IeYwj4CxQCVmPXDGR2K2/0n+EwB8XMP73S0T+ZDdzWb1G8Pnl
srcQBI3E689jZlaxB21PxQuv8xd5fhTgyFde3gi5NwZ9bCD2hMMaOKhlcb+6f0ndBhgCTC/OqJlp
hUsDo+elyX4YyQ/YHb8yaoWN4BpsXfSO34rjtPwUvay4kn5vY1iyQo5U+uRWmZecOWYJDhX1UkcD
TBdR/1XDIqRzAmjYNkgh8YgF9pBNMJ2vxJUxUOe/1p0K0yx50aCrswUteVHHIB2DF9TT10T1Fupy
dZLywtpigxmxnmXrpAqskDCO1Zqt3Knqq6jXHvZd0PCADczHtfXiSXvTP8ZPFtWpCsTUWwQ4THuv
nsxnYyqOno8qeH8BDxexD8t3I+ruIc1hTC6nRPrSXRoKSFBhtBSdKEw4O4oHuwlSfn3hFZby87+m
Z+Twf3agi/gbTSjQRR6AGy/bPwAWjn0C66vMqwsToWSGZHtQp5ihqrqKDiSYdMsKASk5ZoNcpYOO
bt5o9z2KZQhMMapWnGqIq5edv9UXw/M+H12cnzPapCoexxlodRiREOOXWEeiVLItQvZ2KmAQJ1kf
mkCCIxmQzF4LwurwLQR54e8XDGjAfR1QxbXGyMz6/O9k/QsIvvcMCtdxxdFXcUtoCYv69oJyAvsw
MRyzGnPs7okfDGdppPxUgbkGZ5DGewe9mUbyUN6v7dwI12YwRGyi0ZYJddpn4DE00OiyZkIIDs/I
kJdM0MWEzODhN5U+HBuUHBgDOVLH3U0QUCrGASz8FRhJuKP1RvoS2raVs32PMJaV8zdxhJsl2O5i
zfLxSwcB6yo8cOMsKTg0bxV9JLkStT1JJBVsihhrEUX/1e3Bjf1Rjx4ylNkeBQwBye8qYwDmqL/X
1eKK5cuvPEFBi9f/OWdqYoix834ZT/wcuFcsZE/SmC7JXo833d0rmxpuh9JSxpjWkuN3xfInWZJM
0naDlhXoTQPu1kSTyVgWG49ImPEAfYCsC96LJ3By2M889VQ77NuaumnJheBhD/Wf017dlKEBCWxf
3DVO22Xq7jJRtbc5/A6mjmIV1sH1GZhwSHs+0yXn26n9cmAZT5h9s57rsv2RVNb9bThyHN4OQkb0
M+cUqam2BrLM/5wRdN3pVlPQF6dZdyp5M4yQ67D4r9XFhVYS1Cos6VoHYb/1gAN0/PXtV7ST7w0P
DrJMvwwmcuHi4bvhVZdDs3LElbPu/ti1i5RtDdzImaOSNqDvwweFPHPASIh8tFkHxaL3G/VexqWj
Wfv2OpovZ9WtdNVdlx/pzg2xZiDwzajmDJXU/BEJWHAz9u8a3xnPQJLfmpnkg0ohD6r8Dq2JHlH3
MiBJzBimn6PJRR+GF1qbHZ5DCtREm8l9kZDm5SBjXnI0/ocQbyHuImM7ob0UVcy5+MDX60Tmfe4R
6snT0A/WTwGWQfWF9QanLKL2WgqQkmCrvYhedhmuQrBjhY7sNla68Ifm+gb1WbOegbA8NK92Dwco
P9ig70b2gXfqa/Rvv+QBRUEeVLmUJcPJcfRbJdWPr5zR3OtHOr1vV1wzkOFPALnRKIQ69jvUdlWy
hctrAmhqcqSuIIJG0b5OcJt10GcUK+iKlE9quZH41oj75j1Nq5lPc7FXNCM50HC+w1PD135+5o2D
G20eZYAoiEowDRBTJDJBcipUYUUiUW8NlMiONPWm8VTEsZR+zUV4yJMVmJzeUc55pz5u+uR8ToFn
9CMwXclJ8hwT2UpipkLmKPOX+q3SROMriZfcoLqeRd0P3hjnTIyR0Sbn1jHfiTgJXvC39FmUHI77
5ELHyNNnm/RZ9muctJdiUZwjm0Ta0lRRWCZEB6FyQN5eWESd0XCjLA5zvW/CovGCFGijBNT+cDUP
mAWQrCd1z0RlHUgi49go39KoGAX+cWs0c2qidYagLyihKQ15ESrYZ8UTnQEtw7DCgUi2p+CG56Vl
YBdMMfqYxfE+Z54zSSS422djjvbhH1Ln0hrRDnszGp4iu//eKur50FktIiY/WeRlQszlXpMjF8fA
1O4rcFaxQDTFnGAV6t649bmMgC/5573eOuUkwUTa7ovE2rRVM/12n8B7O3Y9PkGzsKXWlKHwvUjb
xnT/+PspgHcIXKkQGtF75BU9YrSiFQNWFOTFMRwKLwUDd3fytHs/jJXWaq+TJuR4AUTeNgSIDBrf
F8hXhhXr7YsfimRaoBKfuP0Tf1yPtqUB9sJv2pRzt/j2doUeyjH3horv6yK554kaZtfc9ae80klv
CGfxa2hpgrfPU7WM1CDut1OmCaNDX3UkPRxzHzJqTe2FXrGZgVvPKaTfnD1sC26OoYPEtuV1DgLQ
pr2IuFp/hleQ7TBCrX+PVn8Y4BkUSHlFTxeAaAPPy3Yw9Iw2vKUMU/61HLO9PvLJRcwa9GryenXC
0CIgHiD1G2XQZteRv11UlUy5LW4wPy7pjWwHkCVO8eBDs18+Jk5/ECz3O1yHpZ5GetHGu82AwSUK
l09aKWVHcVtRoIo/velp+wTVBgMHVchDG/oftkYNI4H4acYrGOqtWdTrw8rMHhiYJct10cBfcrRt
Xa81j7cIXrEzSvltAPXnItO/4VAPgxMPUeeHhH22mqt38KhvJybh8jBhAV0ni9BOkgjs/gqdk1ek
zYmbDtAUw9/EA5lJF0pJhGIlsnDgVPatciJAtpaM3qyPTmxJVoDtTVqu5OVcMxDOS58OW7VOiwMu
nzo/6AYIAaiW+uytB1QY4UnoyryqL5saIIyX8GJ8bS6usLK9Uqsg6Jt8VDymyjmhaPWjptFvZuRO
w8FrrdkbX+TJ69d8cdCW9WHaef1tYEf76To6JJaQ5ZxhMNThFvDjKZhKh7MCxjl2W9J1i3lYNPNp
Jm8MyxXxM354Xi9vIyJgJXEFDAfaSdoGpIsYKaY0hR5pu17m2rjbUO8vz27ZO04D0lFzGgWTmVW9
HUqo1AvfwtjSdJenmbIP7Y+Ebt/MJ1mc9tGkiPn+3Fc7KPkZzs+vh86jetKBE5bnfTiPecacs6th
Z5O4FZ446Y3fYJrUU5YZsWcliCKYseszg+vb5o7qyX761WAPMhSmLJPqAkZeJNkfDitvVH3+tY3D
fBBaoAEELYf7Wm1uuEfINFn18GYnoAJzO7qS/7c9UqA3YopgV3mvvWFtU+KORpJZN19CwHI/vweF
Dc5Vd7A5Zeanv47fWdHIVzFNEwSaZ/TreA2lfpzpPlVFo3ocHlf2NCAuwR7H7x14vlnAI0MgQnND
4tDYTSzULSQVhCTHvrV7loDo3kg+7Ie1aNIblxP0AY6fy1Bg1+y7UVxCCmoYjDtH5fGtXHw3gXxu
lEF3A2mnHw6ER5M/N6e7MLxRxKe8QWvwFVTjw67DCYFbQiYBakbe7FSgSktecj0ncIkKa2nQTcuc
nM8wtH//PHCtDTJy2i+12vtuq1QQeSLgDoo8IHxCkQC80m6p2vJUexpVyVQcZwu79yZpGIJeVGa+
owwo+nQHHKj5lq4pEaC8R3LKAslyBUT+3IFMa2vTMFMrpNFbJZAjTXRJX163vp9/PWVnKLytXZSC
wvWSdP54g6h8FL1nK20Flo2IeCanoKBQ8/m6KO5htMtY+cXatrS1Agdfaw7wRCu98qqDSzfxMeNM
VnoKIgk6WDx2kShcin5i4Abu9DiQMmL5FDO+C/rLlXPZYbGw6BFhiY5TTj7gMFtUeJ4HT5qu9FK5
eb0GXwNnGatbDfO8w+Wdm9XqoUJqa9EVA37uytQ2pYEuWw5E67L2BK+7RdmVvjmBPp9tpftetGe/
UXMe4Ih6nSvuMWzqmZuCVRDarLeDpAI7Jb4gbz6ggzQ0/cYEhFZt9q8vGELQ2GutGZTIXrHlaGcJ
3n+qtUDrETCML9ZrfAtcHmG8mAkWVaf37YnnSGlFWaDX/aXEtb0Y8RdRtwqTeqPDH5uMUOgrCPS8
FUcuWt9tEQQZ39ODTxeeLL7o2I3kmenHC1mUCmDmfW+Q9PgMWosesKM6B9O1Woga+iobenjJ+FPa
rriqYMv+dJwjisMwmla0Wq1j3fDNk2OLvBzoBnNvfJN3d6U44ypOVdU3pU6hyfMlxxz19cQ53O1u
M290aw1Sm77FEYtImVwL4stbNkA32GDC6FYkq3FSdFdrfi4/HTHFsQ6N6oOX51bdySY6G9+WDq73
SxY7Vu5Zf8m9Br93dUmhBKjZmWlHGrITgSC7MnEAcPSKZe3OOaWOgtSz6rpD32g5bER4U6VCdE2q
wrB1E2L3oTN0lKuvObN4j1GGOxFIgSJ45UGjGeRai2joqQ0eku1bVtBT1QbZXOQ0hWSrGOkhUcbG
O3uOICxK1DG9B+6HoMTS3gSOI8thtwNR18iAzW/C79pVCYZKmJZ3ooSH7e9J5Xuj1pwK5dWJLtjW
48rtrq2/Nikr+hHjb69dm0cboTAWnlUZKKLQAnwl777pOtIw3NunKdhVvVRJcv8q3KJFTRxlj8S8
iWi81qtpRcBE3mnZ1xcDv2+0X4Q7yXvwfLPVpGJXJmu3J6ZQ9FfMbR/H/6k+NH//KYkQku2KBko6
vtMTUqKTbJaXu6L9N1zZnIxa28tgzP7JZusFpKwTPNsr6SmrqA56ipf2vxh8ONbYEmwgmOcnkVQs
dJ5/115SrjeRDx1uR4ALz+LTn7m7uxyXFiwg2A67Am+Lt6uccrfY+iVybh1oFy6XM9JWXnYCdJ6D
i0/sUn7/rI5SnPt7pLDaseQAl2V5uryiZANbrpBsRBGQiuuM3hbDLSHHZ5nGiNex3SfUySQLP90R
bMoMmD7B86LTNWn/c+pRqqk+8rPoUTgM5++/x98WbdQXPpc9vxJYVwYdrLd45sVUKbhfdYtTyszx
NwRtZNFwiEAlfmW2MKma2qkj8/4/EhnGIts5PGPVzpdwjFYsjYIONfcQ71Rbsvu9gxfgixSGcQRi
KiYFRU4wF+8Mt38phq4oHQlyb1KEMSvTHmK6b4Bj4ZhSMvIrnZUMaJEAGGVHiF8ovJgxNaSEZyT1
pvG5TWbbXoNo/Js10lY+qFCtGkdztxn8oLdFmjTCARk3YaOjclPfqmPiKglFOWgApJ4CQtTcVgCP
xGBulsZCC4lT0Hz69fGx6ORdIYRt1Ksvc0ubuepL99Fouhl2aTVmLpYHRglGFGJB8AbguP3BlkcN
btBNYepJUfdi2ZYBcHmVVgQCWJkev2JvXh04WEgaN0CgC6cG+sqA/Ih/mtj0+4kH9Wnd7IRDt+WN
yfZDQYSvfuSFf55llmmFUa8HrOCrEq06eKOq+ziE8I++tuicHzNaQHGgApA/6uVivjAUyLvYj09p
AeD1mLCmXOXYRnPwHIGpdxJ2NPU94n0o45M5Rycn1Z+Kl8EyFVfZdAoRaCLyLwaHz8VQkHv77BgI
m66bBFr0GG8n1nKeXCtkBA4zOwVl2ZaxybS4wnYiTwIu3YH5YK1npkPhse5YmAD8ydLEOrO46zYP
YnfmMowUKs0fdKv0vKl8B61dA2LC2HQXX2yzP9Lp44h7JSp3hBINcEESLUu6giqNEy5hGVQTup9b
o0ixCHxBfhiiFXFfk6bXshcYYRD7ma4vfjpNx17psJmuL1X3fGN3TS8TlW4ZboMR0whqxk8gz34b
uviMClkBsG9Ls1InBY/kyErhDaG86ekvgGrB0COnRRDLaiKYHUOzMaEHs2wUjo2Q7LuGQfHvRRSw
wmntFNgJsstvb+p3rKF4jdV9LBkW9ITibwpyD5C7zPx7KpWJAHEbwlIHvndxgou9gvX2GcE306qP
Enuue5+cbdqezVck4lcLuJgdAag2oGjPFmbIzGVB+qfWEcc/SbD5phKjPBgW5YqtXMksinFErwIk
rMhuNUVx8ktmsVXOb7jzlr3PPKnBTNYu38+sYh4W6CqwiyIqXNdzjnJ1YsA/Cx5ZgAtMcGBDOE1J
sg0a9A8wIvb8Op5OuUIsH9hY5Plb3RL+ubCU8VqoQFqVcXlXcE28E7WQ0Aoz7pc49Xa154vakUdu
TC6S7HA3N3h2AQdJf9jXnOjIpOZoulZnhHEDhwKWFzCPEVXyU/TntEO1xT/Qq4g31YraoM5l+2HZ
ZEYSXqKW7e9wKh3d/QJsvfJQVNt53GLt3J3Xp5OWrkDWrC2h7B0Jxc4TX//1/F9ykuEDMcCtJVBK
3fqqGVQORhIisW7ROR+zmk3MORpKzivgDChRe/6Zf5zFqQ+F9UsDzfy2XrTRWRSjeoDykKPD3CT1
d3DNx9bYS5p/IykQgqszwC8tDQ6duKwEFwQp5jERaUB7DMyYVVhWUA1ms2pXHATIr9ek+BfBzSXi
OVcBsJ+bU/vS8eFhxOsIoWLR2tdbaLvPA/Jl72T4kAY4MNh1rvUFk3qDA1OmwxrX6TCuC/lkF2M3
as2eE890KvwR/kKqm1UhdRLiJkEifmSGadyi+ovcCfYoNhvNiigLsqBgEMZrpw9XJtq1413bQw7k
D5NZuz2FgoggcxVBtxyVXUc8wpmJAO3HaMyybvAQmPNgF4UtZ8Gk9sb+staK6GQed1VPDquYIlUd
AWKS0qzcrY0IbxHzL+hpem28G2X9SQfmljAOzWHOW3vYIqSedfclwm8jyY4wkMLwNfJJABMEgJBf
73qOPw/lxm4C2aMpd21eqy3hGe5o8OT/Lgn4M8EvQMFEiafBwW7br6lFsWYjiWnQB4JOqS1moa6t
5Xdwqkb2Y70ynd1YoGxzEqESuNj/IBSYiPSdMDfQuPnibIQLdVPaGTZDQkoVpb1qKYZWEHzLkU5W
8mseAUvHppXYkMEVF/m6GVaeo6S6kFwfKsxREydm+oYn0roQR8C/3NccuH2xba/JA75tHca7Esjc
MnMHXYZuQk63b6Iw49Uejc1LVOqleLcNHFWeLd8qGxv7IGyXd2rC7nUU4ajdzLUUlKgDYLum2dde
ZpUz+gPV2/9LCR4vWm9esCvpojxqIIL4TkCyTeeS7Pg4ZJnHM3GhSFBsyIXCqlX2H3fspiMpJVOS
dnSR/EdI3BHlvDX9PiS5Dee7Rpqcn/GXKbVC8CimX1XGePGM5sRGvtlAu92YJutBuqa3kA+BZCFO
2pMEG3NoVPCxmzvD+8lZkm21ryZXWLpS+zjPCYh50BSO6DXMDWmE1pVXKpM+QnswN+/R+HBmEyy0
9yLze9wPfql8K6BYWcrw28NrDFTb7nVkJfFge+8KDg53bsAQUK5hodLcESXrTdsiVFgQA9/eQ2A1
LTVg8pkuoKAslQXlRsIrpTCATvI3HTqwNb6LXlva7pm1kqoVmySgayjj1p9Jkyxm6o4Cw6o+L9iT
Dg/c39I6U0Lwo+EC4yVeQHE7poywQR3iZeyyz0liROEXIOR21S9C43S4/MnyMLMX7WjhYh9Iym26
TWdsv5Z4zUyBWxQ01ICsETWoh9ciFXkUBHCKa1xibHOw6fy3IFqiXgpPt65kPzebI5XlVb96c23b
TcNB29aTmKMA47lnvZ4Zx69nIo2ijW9Zhv9dLdUv5DqLU8z01GYOj2zFjPMjocXHmnCWpk0sCO02
gv3rnJevq1pyxDUEyH3I7FIVCmqVbw7azZ6QLmsxqfQxpx3nos3cLup8yyZnODTZXll9TYMP1etk
FimetgQWwbFOqUhIf6JrVMKOCMZI6ouWHnvM/w0aGwO/juOhHZeln+v0N5TL4hoDULqtQlFWp0JM
Yd0qDIPrM779+5ZnL+d84lGBEHL2GlP/spEbw16acvySI4kH5UVs2gtAF/Gt7CbSdti8efY6lQnK
S7MH+qun2UPNSCoFmh3SrJrZT/JITicryfRERaqHZ+rDx7bi+1c97QNoOCCeyVdkXofIHkh/31vh
CsH5D8/8dYYKU2bd1xtxEPiXtwTi8pP+FKmcxIuWJJeg+GqlBQlOkACVjT3H8Fw24mkqTcTA+PEC
N5wHBl4foghHnNqRfWGSKmtud9BjubfDu6iFhuvTL+H8gtcZTrappMblmZZWmm0w0hWloqgK+e6j
cldkIfbYdxQiRXpk9fyKs1/i2UsZQt+LvZlZX673cZfXCVaudQEvcLMqOU9nu/S7/Hkzbq4eB/vt
CZNT/Jr4o76v5CfTin2/p+sIVmwhVgBkK+07PdUshj3xMDw3IQn3u1trzPC8VqIlHfptXq1alXUq
jIdH+pHBF0A+06Upw11RQxaZkaMg1m/pevB0QgQau266uf93u481snX3B8PDFYCiVj4bSJIfUBpX
QNnzcwM9hiBTVT/HQuF+9e0c3lwk3TppJkV4JDKTb2lwAYkTQTiBo49LoKBpLayeAx2tskXdgkW7
RXNJTU7Ojii7bZ08Bm7Y45EIpjAmJP2imIZQGC2RzJwcXRduHBszfJXcO7sXm6dsqdM7yWCFVi5m
A2zUWlbxeREGJRbDyMakcPRBRXM1vcMWYVEm9Md+h9t3a7RgZ8qS8DHAaOwzwyVEpMjgqAyP+mf1
2XV3KfD48LY2DGSerNG3Veb2rFicX9wQAJ2CsS2bju7z27ECTRq3X9Dvs4zXxuMNngc3v5Q7fj1i
fqXaSu31VjW1HyY58BfkJMhr+/CO8SnwOSgmW4xwbR4ZzoUXFLXwLh/NCDdb0eRB6vsDu03a8+vV
Z+MGmtBzk/MhaN0Etww4zJBVpLgPryjE6ksOd8BtNcgTYhOmONZO5sPZUvsEpg4dpURg25YE3QWK
01mseNVshPhvNpjFgJ96GL7GWBazls5ReVvwjXEfWKtCFV3pT57+NNd+uVr29RHwubdnU+DegZbl
LRvOtYtohGIue0PrL1ZVdD8jZBwxMLUd3tZ1Dkzm35cO2X0Xl0m5rkKAwDGAwosSiSPlTQ9kv2zB
5r7jCBUdrt/Q/BQdwFM7NjKPpM3xLqu4trKkyyAV0vAuzFjaCdKitJN9ufmncl4VTRRtHxMAJizL
zP9HeOj6youFbTVZK6d4MGvfCeSya1YRkD+IlyTdKtoyvpbiF4Ti1ISEKSd9M47oAUL/8wFnJbNS
4tdkMUFXxyisO4ZuMvzwumak5yykOjqFmDRhrPd3/Gn+lQSgWag13lAxGSkWV2g0iBqRQMprENbQ
9okRZVr0s90ahvfDynI2pqLW87VWF/MjQcCWmX+Y+mHD0e696ucbxAyUY2sbvziQwA3EKvm8jBjA
JZ8TjZKc932JIzllzaZl4Ha+i8CEynWxx2uRxESs/N0YjR2qKgBrwLWK2MHuZz6Ys9x75bbPCi74
lisS/ufScGrvVvSFTVbWDe1gYTGjGJXsZaEXXKDOZkkKikAdz/7SuRrwKDSktGP30Kty3A5yu3tm
z+dCXkLUwwXReZ+s1amkUXJLnrutM9BMZfhQBFe5lpspDWRzXCQEtFKQTwJwZGuBbsiYn6NLB/w9
iab9Xcyk9HSee9U1sBX/pIyec5ooEUBgj+6N6DZRqIQ9dprf+rkOj+so0+mx/TLoHHsobaBkpLry
bnBCCPZM/9rvTip6zkRpwz5b4Eo1g+CfKWJurlsjspBdY/lK6VKYmgdk6TFJ8NXAcFvUaEjCmKaB
d8ptcJqYlUNMQa7+jIjnnHsqd6HfV8DB87c2V3ENd6Efu4K8Si0aQPaJKB/yIOfeePxRAdU7VuvJ
W8qA0r63sAOymFwIRzCQ6L6KRmmOW8MW2pZrStHwL/3Jmo/HjAc1gMfWApl+2CWWhSOCEiKmrcPW
mLf5QR0ml0hZ6Kq/1y1tc8yLKwyVtIIhgFNLruYHCbJXCaqIJT0w7MWi6uuYyzwgXIwlHVMYnv7p
OPDIByzMZp5VIDT+2Qzb28iqOZgmdwxtFk0ZNfmSPEItgIXJpQefabm07JO/vPUdYg2tSYNcY3AC
uAoOm906vVgkaZwEnq1NJhC9B083M0GY8nhZUUyYCAxRxSkGVXmVAen61iCvjBcfl2t4CA08mQGf
Mxaq4ayzBOrF04d18Ofo10kamhhailiV0f/8UlWDb84t+nftZFTQK8hoy5+q4t1HiBjGHYwM0BoX
u9dm1k/GopAvL9MSDTneO4vld4mql2KgJIDYFkA65wt8gAYusSAjXzHhQ65IHt7LDSp2WQxgHG3S
CWKlH0ckKK2ymWeYvgmqf74iOaKab3YiUnRU14qDvGTLnYKrFQQtPsL+eKcjZiALf42b+U+FzX7y
mH8M0UHuimpG4rRKehBPHdrFhYSCnzKf6rNjjt9ZEqEhGcn8xL6F779oFiGPGQHswf+Oi6euCC0N
/yL4DhV2JIszLP9TiOuYG+idzcagaR3hZRV+ohZz5jNhBwP8xSJ7P0jxovH72bJyfMiVahm7tM2k
pY3uVvK1jH00dceee3KcMmGODBlD7vDdM1QYyNsZttN2Lom4MKIdfbht4L2YSNxYbblU/PjvjfFz
p1z98j8rd5RuAVdrodrGI9qGtMdkwM56aAtOqzWX1cDo8H2OpEuPv1SgGQFu9/l2TvWVKo4r6O3m
qXQH4JSTW+TlS7WW9qjxR/Awzk6IiD5gkrm7QGDKOcRxt8cN53uKjwRv0yTV7ddkmqd3g/lDsCON
VcwCxq+1V98iF39sqdu6O01pee36R9ayD/o3uhPaa4d0c00P8r11m3LPBjHI6Z8hKNIY3ZFA11B3
IiT+thmuZlrQUK9+tGzu4iGWJPF+aUoDW6IPzny4yFoMDQy1p6LyHDT940AwF/aa5QFsTIIdm0c9
LhW6+rjE2Ln0bq6y6Tspo6zxh9JEnyLrSgp7HGVJ7qcjO/0pcqXRdSB2XXWsbgKjPmGaibm8HME5
ewhkk5jpozy8eHg3FsaOoBhny5eXG8RW50Eu6fSOOgOPzWTZq+UBDTbG2k2W6H9QtgVScEfpEZsf
2aWIaz+96b3BHglEmIXp7M0pN/JU/R1GuWOQt+bZQgamEmSKhNTrCzobxLuCqL4WwvbOTl5/t9+a
GzduiJafBHJiFv655TNJRlcple7pzWGL64Ze0eOSqT1LEYaodbx8wtR8jTz3u27O3t/folCwNm5z
/osAF7javxmx4cg+rKj7neIbCLOlmuO6KPWdkICq9179d9XcX2Qh+QQHcpNOGhFT5qPMnQ3vR9E8
oqIFUxqw1aC8KV/408Bh5F5Fk7WPXtL/eg7vPZz0ysoVu1Pt8HzNx5GorbJEobAS9Ik8HC+//ko/
8MxiW+SOoat7pSpPqh0LLpUTohZtjWfBu0eMsQSam/obb0vxCU9F2iAqV2dv2dyell0p0YmBkcmE
iIHs5ybSpgacKszZOeCzqBm6FZTrWebHaKPBawAZbHhPvlhPRwrIYGQcCnpff3tTPSdfkFhqbIsV
d0YttTVLsP8NaMKSV4e5AhXiT4QU+I0Eksg7fJ1IWxg6DNlEvkvYAGn/GXCsNPH5j5YLATVSceXj
Eqi1j+/zpI/cL21mB2MvcCMENApCKWulPYsLl1LYzNJlFF9vzWJLfdvuuaild8onTNlihMpjVRQ9
LEa+1zHxXN/JvZwZhjAFFnxrmZPy+3Sj2Jd1Bmje3iNJPBy4eVmlPiWjUYXf/2ZQkOCaBHkCX/DU
gO/tHaqr6Ss78bKTIXEKJWeRrlpCF5KvoA0SKoEr45lAaFvz//6JSbgXqd/E4AKRYZD5wXolwr7P
Qk6J6SQpaecaYPhFkd51xcFaf6yMIT4vPgdfg6NdZYBNEKlX9j5Nb366eyqmpeWbogg0UdoL20Tp
jVPphgCDtq02z4hicaFSm5pK0PenH+qY77jnhQr5WB8PLyk4/naUos2x5UaZHQ2CtAcpu+L9pg2p
DkZA8Hi+bqC304PGxQDQsZtfodSVEKwAZFoW588lmrnUVwlbt9gTjByHtMAoHOBiN7QUkVMrat3K
oXJEmqfMJM9I1MDOHSm+zomsieLje8K6+oAqDSKxaHGbXAtW29E9qTfk5GnT3+0znHT9s7jiuRPU
wRJ1oIillbN8npzULs7OmKCRluP6OacP+SBPFj5Pgmnq3BtuCxFzRcoABzObxtiKYU5o6zLBHlvm
D6Kxg8JPsaasGm3TAb5bMPVOU5F5+kmWPe4oS9DbIEBK97Hjkmt9ZIBq00vn4oEux00VNNhDqR9A
p+JKSrISprNyvb1c2P3WvlyoeSfxPhDSIUdUOtEoBeKoWu3PqRv4pfEBjigysGHdVkafZQrVTS6e
WCGn2BOi7B2qNaSa9TnEDX18tc1skgjON5E8bjIAF0T9D46YVGowGArG8nfammucC9mtqWiGnDPq
EoDevvrWNsnvgnx6St20NGPDsBv7Y3xVbOxiQmUbeMpqF2Fm62rJrV7Zw3IhKn0ISzS5s34avxxU
/RDodjLVZ98GfkH9IUuNzcvkk5MFoCN6SozIFqeZzWvSPgbzdrNrcOs0qFb+O9Ay/XuHBG71L1LR
cvtymkf1f7gIfbgJPUImtqSD5OAX8Hoq+nU0F3CqVC9Yjr9GE9IqwPO+J2eayiYHGj0ucECwsbkS
rU6fPXGHKlWPl8H+r7QAuIfywYcV33vwCwabM7jP2I9ZahNrO6QBwUmrxEWIWcDc62yaC6/HcLQF
Lcz9Zy6INWbvRUEVBg2hB9oPufbUk/PTygB2Tp7dPORzWWAMgsFwoRcVXxNyx8QY+etIfXiew9lN
2Ez3YF2rMyBLduVOxO5E/RNzrh9ICHNyifYkUA1XsuKHnvCFIgsYHOKxtU00rTjtSLCobhOyoCDR
MGkLDK6EcZBOahZTaimBNXF0i8Ravtpp2dgrZ/jdEf6s/Yn96dEMot7GsoeHAR+3pDpFQRr0+g+J
8jFBXrtXwu+pI/aE8BG3sGrLAfwAOZ8F1aM6ozNqPqweb5DuNgbjwciR8HUVzGJSkpWavdzHjscW
3WfM+gLQXA45Z6mDoJWHDQuUYZAomqBr1Bc3NxlC7JOVQffIsjFgZDyHdTWFkZ0YUniukKMxxwzV
CCrz/Xa0gbPQwAaeHSTuk1D5VgfGPsGj7eiUnQDr0XKsEdHKMWnRiowua7N80fbYEpgiYNJNHYeA
WUIs4U4vp/dlw8caAKqCq8146hOM5INV9ju61isqCntrpI9SjTVki8x6osKlCfnmjxZtvlMJm5pg
zeNXnIxaof8V9fpRf3oz/qYbfB+3FR7kEqUuSvGG6JZ/iNULvF6WHOVKeGQOMlAKcOlg5x98al/o
2TgLjl/Lt3O7CZELHKRRRnsL8aZnyTKhPhJD33DoiOj+9VLYSFeMWL+vP1Ph74EJUGB83Mw8YV3D
mqlVgeQvalIn/YD+iDZj1ksPS8J6SnqcYRo4qEd3o1Mo2PjTh8WWiCE8LFJPR4Tf/jHDaEq2eRZ9
RfKVmntTz9+Cd6O1LxZZ8DR6Zm8SIp5GtWnXZHz3TTJie3v2TTDrENSqqxiAVd2EkTC4sNknDgwE
0QCAUmNR4fUE/DLAX8x5kKnIOBLPxatOtQK9lyBqgTBa8BSQDTH7XKoOTK+k0EL7UAiTJ9bceOwW
tLif4zlPxzDhipV0yVYEciogYYTDiUNOw05f8qOfG+zFHC8x9V60Z7Wz3ArFF/CSOm6zuzy/wIVu
5pqvgwR7uISqS5J8BGF1tKIpyJnsbGTt0tEjFy/brRhxMhB3syOb7z7ZyCNbkFJ+DAl3SsK6HR6p
YlLjWiSxIk3ENDYIRmGdGQW0KWquwWxGCZFfTS6giy4mUixZLmdQVJt31G80RIlNhSZ2RYA+QQkj
brNh/JTb7wPKVRTkw+z9C1dCYRmQ17yDqwWN8ADKBe1UectnSrczSdmWdQ4eeGjS6QOsHAhgxAw9
Q6USKpqTRMmTScHrEfWVG3YvcOg/wMP4HK050UcHvQUK/5I278XT4OvqAF8CRfweDuzpGAlKcjSd
BT1JWNHP+DTUPRWiDbSpNarmsoM7Mr0cq8ATO2bgaJgnII8HtV8CpIUDwZiqNfW6IuGpU+E4gYrj
gEXDPvVqQ7uaLxVigAYbKDxRlbUAwaB/oAHEaOiJzpdGNCmFkdgwg9UnKC6hLAISWBCEnpjzJfwk
yFjQiko80NvvjgoQx3EIfW5tTBU6xmVL5I5bGx2VL1uUUHVNfY0SI1L7xmDstas1yMS8NzPDZXWx
Tw6KbHc0pA7CthBkmDRsDJ+a0OQqRobrnYDporpY3Ri4X/BDa8yUPie3lT8DNed9OO46EewkFxLz
sGBTMDKDCxrJcSYCL12i9pdcZgzPTCMKcdKeFwBOJ6DGjPFEePXt53DzJ7Ms/4sjSOTH5SEJsWDv
wec191xaxjHAEDTVzhJEt9LjRqtt41SsPF5Skw4WR8uRFPO9pJfIMCKdftYwjkdTgFqWxvHsM+QZ
2CEzS16IVWRWXhlQst+8WiHsvA7rSDQ0qNRFxY/U64PF2jcz7Jz8WKaW/uAX2cBfmkMUOillOiK4
fE4K0gZZRQ5YXcJ807yXGzF5pSIKK+zh6kc4+DMmzyH0zgI67lTLNzUtwBERac4P6VH8Qbn7VHqL
jotI9HM9balgxz0DhGMmd8d76cXQ0jKxK3zXuPXt3cLvYRkcHg3gfnhpCO3sk14OM1xojG6IT7Qf
cza5ZLd9rkUxyFFL0GpyLln345t8eO0f2seXMDaPL0oOC8SaFNZxEIqDJIkKTEwx8VUKZDS6FMYe
4jVbok0ml3sh+b3wkhowoVL4dk0Gz4UMZdjkKQI6xVAKIaDYdikMjMB3nFIv8IDiIv2gqtCwgIKB
xQ6W6SvDXum1ODSXqSL1fdCOdiRuypd/gKcXTTpEDRRqdXU+hZsA2Wyf43mDcbgS/wNw0F+VYd8Z
6wexVGUEf1ibawEA0SrzXsKHEo7r7TaZ/Gh+ryq/hEVhKx36OGKy78RfBxsOYD7U3d+rpEVtAL3F
OVOQP84zDuCCH7/qxYK4oiMC2BqNmahyh9Ktoaxur1D7k4sg/fS3u4wgbCg3KuxvXlJkXFxW2Boz
D1UWMO2wZTDomzoI9VrlKmkQWV/ORtNUKYi4s27g4fkGbCcQHp+jxbjBrMMdWcSNXR9ytXsjGUsM
FJYjIh9TH5UV4m0s2VxBVShUp3BKEEzed6emXbhnW6ToXEeI5eS9UDRv/bC35jvoNkX5IObJu/Xl
3e6PN3mdv8XYrLb4/ODk2bp+XgRdXvFMqsHHd8881ML9GzToY53s6/CAcR3W/GO4FdycEU3TIy2r
c7ES80h8jxksvfgbkH7xgJOFiMlwt1QrNf63wjjAEUUipsqkQkkodlp3yhc9t/dQ+DZUEnsRg79Z
xeTde+Fh6htK7kquY9xOv9PWHKEoR+N2qiZjO5yLnDJ7w9lqBT0N3PwuhYftOdTeQOIO2pH/R96G
Ls7JYMOtLvUDOHAvVaS/c/s7NABL0PYAxk5ASLV/8eEgYV9V/i/zjVtujLzK04BEn6ZbZF4Qdz7r
ih7KzWxUMODBTAn2I6d8OLzfPvZKP3QAXlP3qK7ELrf7XXPFMLQn5xxQ58So+dXLWGXY9E9dvFsD
QrokY55ziH2QZIIujHh3hlSNGGijFYB7Gg4sgkYRnVC8qP72rL2Rq0xPAw1NvMWbaupE+6cigD8F
pvL0UrD7jNYEjNuuTZgIkX199Jm+SMGlemvw1lrw6Hw2YpLVagoZBZOS18sefW1iyc/payzQzI5e
22pskP4SULk3QUUCOq+ctx8otLW4GR9Ox8Rl5y+0Jj892uLHutKu0GVxe/FfrhtElXhf+pIq7vsy
UvT9JfmaEP3q8ohKjKsjVeqj0GsKvarwFxJbhNApuq/8nmczM+Ow99CDcLgZ33e2vdUV4enl4LFa
I1XrjgIu+T0pmAZPgVXhFK1nfby0ecLXauF8/zFAs/hCMTCY1KZQEF+QC+9g0cdCSNcTcu3Lqz9g
bzOXnv+4OMCXylp7iQf/ckF+5AFXmAPm+iVAbLSUlUq5QnOY8SYCSxw+Ozgb3K6Kjxt54+fzVfHx
BPfkZfReSMh38o24FuuAnBT8xMSNPc4BMG5DpvrdVRUxYL9yAF76IG1Yk5WugxeOIg0obwdjQUCh
E+bEfrWHbFFHaYEdV87iHqdkmEYrvCz5jtNdH7NSp3RchILXF0Zi6lVzxSUL2N9e1GVBNjNKZDXo
oGY7KgKD3IJrfqlh5CXk0ZmcddtlRj82MCfkAAa7d3Bes6TzvOWHOHRSaaJ3ZN3KbyJoOTzvocZ1
hF2dEfrqiEDOCaMGzAtHwWWBS5og7wZOUA93/cETZO/PPz+cdFS86/PuV+TAiNnCRQqMhXrsv/Ro
4LhVzzi8eoSq5O87DEmgEMYGl7Fw4k3Ki8hKG1MxiIVbz06UuKnBnccA73GeHsZ92VU27GMEiIZp
bLn79Ns6l4UVVfV3585sBqge1YWkMPur9ckO4nfknrosSwZa/nCcSGqa31CyHuh6Jw8o5wVLT4B1
eCMjc7ihv7QdpkSTww9pAxeh8Ocp/XyaM/ogfYCR7rgQ87sKDUwxnz5i24AzpEzCx+UCVAMDMNcn
quiMBo0nts4QYjqt+exy6kSCHI6moBHYaVvRHoHsV5V6XsGuZ3ZVYkdzxbWOjQFUMDeKignLqaIv
gbnvZEeCZQK2wtFaDYgqi8L7Q6ih8aVAM59UKkkZTR4caSO22sDSO6YosgYX5949f1Z+MWWbC7zo
tDriKC+eXQyRFd0on2wVOcmtjXev6cgwdEHV3b8XblTWwKzjC8F+5i8BcokVE3t8HyazVTeaoZmZ
QS1PL2fVt7c3PhWsYtbua3TmVVVcHt/mcmEn5EejWiGMjlOq3eOtBObyDrlylNiEG7wCV4WJQ5jr
gZXzWJ6siwp/AUVBBfddKDU0h/+G+pyq3RhtXKv1Er+lyAQxuqlDhPbrKPq4IZw19s90J0s7PVWm
p+6/Mn1++sEJK16NhrvdL23x+6NNW/RsOW/MC/jEr79Xa5OPQgj3ifvjAwEB95SxO82V/ABb+EJd
L29TE88RATfHKTECidSjVaxCBEXef/hao3nXAQ/Ro+YMvvh20rN/aR2S20TT0h7Q24tz/leqzL7D
au0fOLmzxsXaXw8mGo58Jq2rdttgd0TuLnB/Cp2+f3a8/3RIIBB6Hkf6xehH+X8B9/UEbYvBZIVf
YPnkDK2OYg9/QOHpDwldD27S6UtnfMHjNuskPW1429W2rONbi4zo9xYNW8ViKdPGP8LWhEGMsExr
w2FLly5U2epExCcfQWFlcxanmCLKdkUdyFN1Kcl8A2kuySF/2yPi0ZFSo2lHSZKURQG8EeQ1SlK7
XPWFHqZq1WlvD8wLQYyV+E3VULDjhfs1sXHWVZW2Ae/jP8rwlMpg39b6PGZvY8MAxLYBh+GdZbk9
8qRcmPZucfPEtxdG0sCg8tE6080+1xO/aZ3JoZGL1T+wSClAEMiq15IApoWMOGWIIQX7BhueZK18
s5nlDqCz0AbhukZt5lRXEWw0G9k1dtggHzCqUNDxlkGo6H6trrUsTQDQIDHfoijCY5BDdf94X0Iv
Yrp074irBgDV0CBRJ2caKkoamxB76EhXt86X/YafysBFKm83k6jFgasP9EqhiiAHiP7UmnTJguR0
qTjSpufmu55EuTGAZoAqn0jRi+jURp81xImJIz9iGnOlbWNpLfLPIdOvquE6o+VpqKUiIaTCRVYY
Y9/Ivn0EC60aHPBUWhy0f2LnZKby0Hot4/BwU3Ndsvwpwr7rGnOY6fnEg2syNECi6d0Oa1bFMnqr
kI93TAZiT9JWoG2LIGtcDyKN8VSyv7fVCOmCZyirZly29FdQln/7hnJ3GsvFbeV+/W8g57sqaqFs
QIZXZ99Ftywf8hrS7AtDbOirJDWlEDIzG1C4VIH2zQ6SMvXW+7NxZaLB6bO6nINGmzuOdyULNwk2
jRXoHHbNss2IBDKuToOtpYt9jjO8K85g3x9g2639LAVcgrEENlPcklxWVBm8XOaKD9z4KoBHIW8M
gufmPLivp2lt4rf4NdrJBwpFGyfJ3LTnViDrD/pkCwTjznkSaBp2tt4uez3r398P/YOqfgNcx9hk
6tYh9g5Xwl/lGTVG95wqbyjorO0PW7oZ/xjuOY9b+gtfa4TEC2lZZXE8i2IroXcn+drroSqXxwME
lnM0Wm0YbEfO2U7sYDMbLWUXfInsdY9UNkXGyulf4ev2fXI/gtrWcgmFEVHM5tHXotpg9MOf+Wt6
451YZ/oWM2X7S9rglzigbe/UG/V95bmDQ4iJzoIgHWhgv/9pfUM77r+WHQdzAh3m+rJxDumT5sX0
OTWuYDbX3NkB7FELd6W4Oa69ThuZu7pO3Xx0FMhpUtskIknJRQgHRjEoojHlA+qTKOasjtLZNlzL
2oOdJ2dCsVvxLtpr2PQFg5J2cSJ29CYapkKBw4IrCBq+bSn+DvoNR21P3Q4SMSe7widu8J9zNi39
u1OKsDiBxeA1v10dm/lzPDPdd/SIh/tWif1WcEXM1stF0Sk8alP+FVo5nYulqErgRR/7hCxsh5mT
uSg4BshX9yRYpYhTiniy4XDl22Jmk5wlKe2/IHwfUQXLap4dYqE5iNscGvsbU4pmQkUuruiSqZrm
e3xCqbBrr/rUszJbPe6noT5G5Egh9OKi4BnBvgjPoDeppIUuX1+uFxuPi2RmcGAkX1I1sKf7vNtz
pBcfXrE7Ly39JFA5g/ribNu/6ofDUL95kwjPmok8Tsazcxr8cTro2rYXLDSku0igbIQ7h2r7hAt4
/NLNexT/alekR3VQBhfcvtuTaA9zFY4cA/RH4FGrgS1j3q6TVBe2UjtGadA2TDfpLEZ3nc7ftp7M
raW/l+m6gtK58+q0wdmSp5GfQ/LHEHCHSQy8soAJ5gsKbbuxusRS1FkalQZfuGByzP3pjR8g6l8W
Te/89R/ZltFPlns7/1YfR1MZRS0/eWyoatMU7OyUUb7obccn3kVzctrGY00a8aF86LnoTx1w/ck1
q+JqhTC7gtYUV1MWaneVTf74h6XCnJ30wcnOA0tsViD+CFizjwA7tVe5CDG0xytcdaNBlGmmBFG6
pXoDwiqw6Hg5KqdTdxuMP8TTny+ENvbvh1KEBwupPd63K3haGKJQXZQi7BAG6ZWQ+7mWgMtRh2XB
1Z+1FauzX3ayJRUSrmOgruNGsuJLn+sJzRR5SQ03Vfpx5OtwS2t5oZo90uWxF2xvKwW9zFCcUlXZ
v8miWM4hkYGMEMcwvkmO3ELcMqKaOY5JPCmOc4hWAJCPnkTO/f5zIIWE3yv6YiAKZ3XS/JRdj1p1
IS+qCP20VTnBgOlHRIr2eZPb/108v1NWHIr/+sG/YlBEPlWtsnB1VSnUc186moy0h5eVqH8x+8x6
cFyVk7pOdO7FNrg4In2wdfo1Iug66WcVjg/u3K3IgAENjzRKfLRa4+Ktk4H8uM6yOmSM2/Ljr7+2
0tV7n1SjADTs1FA00tDjvZHNyaC2MsyT+Z/lSVmsNkXNkexoe4i7JiPCossiHln7lcOflQOvJc++
qf63N3eB1CD+dN4lkPlv4KiMscp5T9CRXY/QheuuvaK3fNyN0YY1NXWEhvnnSGmzYXaVhVZTsfi/
pZ9tGY6yJh//ftu9gGT7LSOYqdAMuQkCqbTEX/fc30jdx2AQembDyLlKkzojbnt04eKxwr9Kk1DY
ey7FwDl0gDrQayjzn46aPKSOvpINUWOgpdv7DPOgsupLSkUxX/4ymXTyBWscclVuGD2/ZqTr3wo2
y8HJrSgALTb1sTGp595SKEIyKfJx34hyUC6W/WKiiAkuKogqWa2HTDYXFZIX8xG0nI4mcBFuy810
q555nhwGv/Gx3Ximp34MMscu/WYYOxOX6eGmsVMV7ybblrhI95pb7/Hlu4/KTur3Y4YcyzSRpFqr
sqUm9MIUviVN/rReLzfuqYDrGtWiiSlo0FKtPHD5Hm9OEUUnOH2Zv1BEamqwbnD9x8mvJoOSluJ+
FkaAQb7s6XdcAkoj+YUUjtFDu4iBOW6xT0X6OjpInOscXpua+Mju8A84JhuUbMg+3KqGuno97c24
QFFVsaY+JGWcqmZi4pBtAw9nUPkBOtFTiIXxGaAwgchgcfI0XnzuOmbwKT/o/iQLxAd4QvcSR8cR
Ng/BjL5zq/G1syFGAMnXiif/U/N0WOcA1zr3CCWDW+MSxopi0IeQ12oPwxJxmVLpmxnszMGO8n4K
llmzEWVduw9FOAISZ1+dmXHhjcaFQuVBMFLPHBDdCUGiYWqgicr8/1nKrSSgUniTgTxpB2aPByEj
pTyE3CzSkVJNtS396bQWtqyF1gcYfGeXM0Vg6qDsRpQOs8s1LgAtkrS+WN8fpUdKGHfR5avLOhkN
kTgRZ5PA3nfJxQyYa0xIlvmoON/NTs8LXIDx7st2Ea/A8T8MvPNrEGzid7td8IL1x9batDo6I9cY
z95a1IQKUwkqyP/gvv5TdIXDf7ufgtYA/VT/eckBNBA8WHxildJXS72e1WWdWpI1LHhxENVXo/v/
N1RFxTUmUVk5ravTR7fr9rVZp8IhC46gOo3hDsqufkT5lBq9gEZDwevAyucZ2S6CBKq1yTn7og+S
q95/Vd1sZyJi7X2lFJOf6bhxW6E0f5Ue0gx1B4daFh5FChFodnVkEl5ruge5QUwDFH/xKsmV/Jfj
VmbMhotM64oKgZ2vxJRRctdoeY0+h+thOWzgxQHX1X4vlQIY4nNXrCkKq//u9Xrj57VFmwG216du
HWwHgc7+c/Hz1UyUtUmAueW+mLtS0IKSYI/CAfZuQ6n4JWiMaGAVOwu8uFrkGHpRDmfl3fyt7CbR
NmjJSoZ7H+XlqxQE/qG/lXoRmwjj6IthxW5w9/3L/vS+ZfgkuQV28Sc6QWX6mSgzHm5qGxRHRAL3
8YpmKDBbxPLeCt/2+lteK+EUvqgfQvs5pPyur0O0VOUOEKeil5pZe5DjUgDQs4SZAJqbmSDc+qOC
R2sHfzx28ulGQJ3IpBEmPTsw3mjhS6eiNIRBDHh2x1GzyAG+l8uXo7xZiVfocE9tFtoFdCrrmP8m
AXlGFHSfgxdly3vykWwMc+2XBGcf0U/f/ScsbtcfgjlGu/U59U16PjYKPx6cn5F8Kca2fSbTGSJA
eYDjtKRVfO/4hC3YEB3apmzaz8Gij1V3+ThZpjCP4/uftnQXZxdiPJYqwDQHlvLgGa2UDEWRIIRI
QLS37pz5a6tUzNrOC2p6BUT2/8We5zzaqWCeqO+Zkbr0BA0l5OevRm9Wm7KiiROHZCHR0jbw1wxI
VtYbbS90pIWe0NAmM2vFk0wji2JvavTutHey5oZMq3+SWNsjZqoDOuH1GH2HK2Rh11ecUjYBM0Nn
t1b+lt9KbVuTMwH1xgply1tyQsD9eKvNYxpsVQ9eo43dYYssYRXsaCuf2fD/pNERMR9H2iqPGCzh
XJ24y00Sdced/8DkqM4GwNn+5IVRhwEpW9SGenE0Q2o9PynwMUHazIH9z3N9DyHy5rv9IjDXfprR
HzygUE1PKwdJOGtDvN//2uhuvtdeOyRDkJMXHmRtDxJc8n8YUFhWZvHhtlhJmrh4ibysnyZ/D7i5
7pK2YRB/BUI342RVsNhhoPbIN3/TII6Ce8uNGpCJrsqxpduXUphllnHJVH5kmu8p8HJ63DOvVe7+
gXeYV0lRCrXKjdxuqAy38bNObwnsmLpqpAWvPvBE3+7zZmkMetzjEsjwjD1rLvSKOCjOGtDsCW/5
cNNbBE6Oi9dPlQsuSrNFDYAWKIMd9mwsPgtE13KtDS2o56AKIFb/H/Fc7JKWtt3ixE4HAjG8tCxi
FIT5Reo4mqRVkn+GsEmHAaTStF2QVUKWrLkgM/62NE3VY4OTsVj1IqURv02dYipJQX8H42os9p6l
ik+ac9R3e4QP2XWZ5VCtoWVs8yeWn6XwwEjGFF4IBzUODDP72gjdRnQkfY3k/+G7NIywa2HuJayE
bbLoCTKKsJuJagKoNcjyhGdMu1K5mzOpI7Cqjtu8FxBwbgugW03qonvUpGwPBDVqNvvrSbu1SJFS
mRisGvpER90VuE93OTl66l75BjoFslVwESR4wJElCE4Q1Vm0afVL83hg7sFA4FF2okqQ4Lx5a6/f
EHKgiqw7QHIdk/w692u4gv5bYo4FDaE02a7Q+jyoLfrCNX/os+y5cA6hewhFfkMCyZ5Qu47DzncS
06bDk5xZt1+gw8Pe9XBheinL67ooDq0S+hq5GZRVTbW3BsOUqoWCXf58hBUzcgeOA0jDkLpPkBRf
gux8XAGI5Ms8RxEfAiulWmr3xGgn2yp5Yhj/P2PtEi8+Oi+wFb3s0ZIeqKRDfa1Iq2KD4KpErxwG
PPwXGSfiR2ofPTswZxwSPYwF3tN9X0hnGlYBaYdRaaT1aTe0to/wf+9VdkzZptdtnRCmiMe2TqCg
eiMUFTvro2owdgYx8cUOC3qI2i1xCxa/JS7pDBxofGoB44h6zqyyArUFXF1dB5TF9UOyGqPBtAne
L6EZmR3uvnNzx5OKNgEDWB2xeEm60Lf9BQk/kuU9LvmUEDhq+d1BHPXFYfEfRYdNqJJ85/OBum28
Q8oJi0A0n/U6QP643rF5YsKsuwGagJZXN1WTU0renoPKwzH4NKlK90C5sQFqPjEwGHUY6w4MrsGf
58fKPdBPrsB6wp3iNziwIamQsaklBKr8rgBNrMxhUUdp7AMcsnD4z/YIw78lg/xJ4oD8UDiCrGrl
kLvc8EVwt/qsn7TkQCyQpQ2TWwcFbYyz+sz5NkIIi/DXpPKPItP+8eh0Qgb3XE31ndEX+yb53jZI
WbbGNc6ewrU6EpZAYebuhMxXPBGiGh3Lb8FCD+jkc8vskwZyGN06gg5xKLnvALwYXfnRUbHHfS2Z
9sGB7Okd6fna5c8+g1P6UNMHK2Zqc0rNSc4T2jDXfRY6VyaAujOhH2fk1YmcqhGh/IzV5IUUz1H0
O8cIYxGmabZIRS9IA6Se0XJqxu2wCSC3eW/ZuY0LQ9KToRoGGLwu4m3c6YKfU3KfNAJ9Yr8Pw+7j
2CHLcdSOCkQ4fV4r/vSozWQwAPzcK0hvi6GNel70piAhEGBvVb7/uAeoi4S4D4iGmg55JqpirBEH
lfx7rvwekkduc5CfMWpE2IGvs3hE7MWlqctDPDN1GnWsFOSyMT4LurRn61P/XdmU1XeRR+r89lc8
LTf0lXnsFYLq2zqJU4+fE1uUaxTi87YhZRhLPmO4R4gUndnDYfy4rQtsEogJPGbYN8v9OCJxUc1H
1Bi5sIWIpU1bNmcn4QB8bZ09NpgUoF/pIOCAG57Ssk7hgC+4iQQKDqiMCyO0qD3lGZLabdNsXoGl
MTViMcxrV1ipyAPMYQxnrusvFJudn3zjUepCWoI+X+5GpS0mV2ADKC8Wxnis63Ph7/cQX57rRunq
bdYm/2JlaLsLPa+rpuAcZ+69E5ytEl7SoGW76FOJ6hCMvL197tkCfpC8a0Gj3Qi8TMAw7HMkojaJ
O9j20JTEY8+8zO2ZhidVM/E9JKhU/cFYuM18vAQB3AodHKeI25Mia9rKYoqzFbu1beMSBH9O3E1n
9RLo/HlY81tpSOCkqqu9j8DITnKL6U+4UynDdf/tyyZVGWsy+AyVlpbxfKZjjq9ivjWilokMJHSC
BfMZ6XblHFdYd5dHvRUU24sWWf0I76fQjloTdZlWN4/BG1gxmYuRyHisLw+m4occfuJpSc3EghJq
SoZMkAv/lIXBU0adFYNJaZJV8McI0Z6HS0uPjgB75z8NzMWW1Pd/iMAC0Tw0jVdOIow0ujxiH7XU
vw+CG3TAzW+ighFoIcQjOBIgJnHJhBNycWFTy+1RwP9ug/I/7vyoqGzD8ZkfFQzFZwXtpea84IKU
KSowaHjULtEh2UXHRrOu8DV5ngd3bSrfoDd+jvogWZ19nOSXuUgCrXAoS/Tyi2DnimsV4Z1EnLvE
gaJHG1g1DfCR9l3jbWtIwrbEl4xQHz2wvcNbcmveFAFq9Ta1/fB7/Ix2eKacMLBtImGoRfaJjABA
U23tU1eKn33spBUAsIvY60Jvjv83w+T/ZCwTqSmpBQE2dJlZv6O+J+nOtas6cUxPS3xzOrHuxWB0
L/QepfatWoRdV/BsTFxNTzn+nDIkiN6lB/AM1+zsOF5h+Bii5hIM1ZbfIDBkMWNNH9RSKTNxJGTS
YKRFsFkevk31qcCd2wn9UOvI06tYOmXKDhFuVllNDd06Dg3Eb9G8CcLot4PWLNQsnqPhQTUc/g8w
n1aGRmfAVhqA6U11VYYLkxUi45hiY85aoxm0dRAyczoZpnhiD6eQC2eCAemNfFTz7N2RLFYXF2fj
loicn7ZyZ8T/eWX+gunPABIVgPaJ+ZMj8+TPGeTr6MJaRBbI0efIFerJSa8p7cVkJiG4OOhN2gZY
wuAJY1TfXn1mPDUgE77u5uezoI8O5VrOq46HoIM2Z8bhVNgBtOPl+jPKBuwvS19T9ZdhzT/jjJgC
B+P+lDKtKoC2VGaMB701fy3sM0+kFUr2HRHkfU4uuuqGtFyZwbqDTjn5dc8OHvGWDIBujyQH8l55
OPSIcnA5UC4X3K2DxXo/gqIgokujr50TTEBM0BciFaH2LfvzxzOkVZGJa9Ma0J13r9O3+gGgOQW5
aROwp3sx8Kw/oj66Wep7nPs0UDorU4qeKsD4cCirjQ7KKmyEQSZzqqevsj9qPBkmJjrwuhKN7w/J
xMKkRhe0omjS7o/Waqjn5V0kUVGsmgmnezN6GJihG/QFYWLCLV1ixOTlAP+Ls747XvsKnS0rdN9u
hQLck285ka9hdbp4zkGwU5wuo427VOrJHQo+sDhOiiec/8lG/w72PwqGRy5IvAzzC1PH/psSeS+O
TceXMFF7OMi/DvsMfYEcmQI08WrrdACgk4pkdC3hsTNZ+lafaIdJPBn7NJVAkDR3layJ9MLB9ddv
3fJ3zMa5L8ZEQjL9c/HbQfGjIg9TAAESiIt0TGhmNGewV7mmeUdM2ZD3eP/Nj5pdU78tneHXv79L
2KWDnBQSQouKrM5Jv7iMPJqjSfwzl3JSM6FfFgMmEuOv2ycuBZh7DmeQYYBd0ndII2BkpxNxZ6n/
4bukeJfZ4bg+HXV1rhnfForK418GX6XibiqHKHaBMOhIBqtNHQ04pDMQcpPXD7aoWi1j+3sjChfi
hLL/d1y6YJAAYNl0ZAQBvCse+sxB2rAPeH/I1QDPrwm5IfzHmIM8Dokq9929F7DM9i2Iv6eY0aUC
DXg4TTuvAGrMc3dL8qhgLj1H/rcoqU7ff25hzVX3uMU7Wj80yOlBIc6xYanbtOdodeJkCFC6bghd
jWzLHaVH0CANPGRka0eYSz5lo1PV1fzcOKfdHscYawEk7S6iEaFku1IutGpL4BBir8JR+juDiya1
hym8eGPbZENvesEQoox8SAPgzV0HplS7EBrtLepoCB+pjH4LnZdX426E31BHQiG7bfyD8bXu+ZOz
vP/zmT3M7o5xNpNtbDn34fLYHO5P+/W1r0zFc534Z/FdT9I5Dis08z7X8eJjJk6yOL6Mdui3rjw7
9sbO7f3iBmiwGhWsNqqTDEBUc6hvKW/rMLJIcU9Mcg9QU3w3T0Gwmk9i/uyromQkcQe+s5zPtw9n
CuLKt2fFWxcm+zbf4tbCXgmrUhQ6Xxu/+LJf711NnXGI7QBT5GQyhUw+WwvGO1LIKI/EH5kW9RaA
DVQX063NWv/X/qxQeyBEWnEUMpMOheknZrdJS1fI6nxTXEwgygPKeISjjkquvRPgEJ47d5jByahH
+LSjH6xZgcsFaKg/0Wmx66oDaUp7IYeO+OQ1qQmy3320fKp5L+5OOBgpxoQl3fPnptOELT7ZkamU
oKV9j9Q9myfnabTPoGS9AH/NMr7nOK++VpNtoU4YWVnD8VUv2UbWp2+jmCRgnM94oB6D4vHzH4HS
BAU/UK8sgujFgiIp9kVYvx6M9RuRdJMTuKXaefMAy8kh9UHzUWvj5s+iPZ9FE8weF13BZlFEjk3T
CffN7SSSJrDW9wG6wFSCVR/JHoy37YFjt/VYO2j/k1Uk0VAU5ADZTLAoaF1fv9afA+zadFhJU0aL
LKKVMPzee7AX49fFwy4unG8bgv52znurQwUxw4mD7pDVhVOSECr+XjExr3ghViXJqyEddhlqXo7R
NkquGLDIroiAmeEFIpKBtgGq794ZK5yFeNPJcLSFSLDnvLYozFtvAOC67DCklnWZ9jlOzbzE+p1y
VRVfnCTbh4Bv3I/r7ZZcLkTg9MUidLXvUeRjftmoh6i30nsv5ZPPhlguBIhK7tZVQE7ALzx2X2by
Z0JrHLVv+WcjcmgQRwssz5CwdJEDEqnNUl5mMERtWVz3RASuCe/m7uN+/0bxWJvsYMgpCBsLhhpR
jnHDoDyoooS2q1NJBIsu3HXx1Ru0b+zyw6PmMEaUMAAJ5VaB6t/IqhaZ7+7pb1vUXNZ+QmlgZo8v
0NHYbXZ5i9EIy7CttWnILy/Xgy92TwYOoVMvHfk3whoRybD5Ubq64w6nvBGCijRG8Rs2/yT60fCT
rIrP+OWARqoR6C937XNuZ9skAyrlUGX/bbJd3RawhcZKtLWZnLaLYKiW3ldDgd+xXvKcGaLRYSVf
VwXFN7Cs5gQ6cEHaddv4RtL9IwpBls81J4iqVdgxYi/zLT/6iZDqnviPoOlYYY5A/B72/RtvLIvE
RwooTkie3d55e5JGUqbzIbpWQ6tPKntAlFU+zK7e40Awo85x8AL+wtUMbftb7KHknsnHMBwVkVeD
wdN5w2UtKodkwrYAOSlyyGwdS9rLHjkKCDvZNVnB6dqdMZO9jWMIML7xhnepIwY4nrDgXYS644+J
x/b4IVBrHAhgy8d+fG9qW8ClY12x2sZpcWXigAFPuBveV7f4adIcSHW6ezuzj7lS+8Je/3zmIbNa
tkr3eT5PmW1GBoKk/gpp3wsOk2cFIJ4UNo9Gd9qzsAScMphs5edGmQKtEhZiV13FXknc0XuC1slG
qts2Ey/HLYY76HOJ9zI8Q/DggVS91t+LDiJHUmR9xzpde2lp2V0nf88f6CJfRzjaouZSnXorT3zA
NtomjWhfQEX+PC1mGj0avXniUGh8lqFo/Jez4pXFcFGi4WzDS6U44V6UZKTby7uAHAaFxQ0K5tcy
Ig99s2ZU7cxpvBZXUzz8dF2MkOBJlOGnk5smGMidJ1A2hQovVHYwzepW3EYpkrdX28sZ38xzcxHI
LDCugPOYF1+plWG7VdVChiqA8gRuqFYQkSJ2IYZuuHNZ5Sxiotx8HvrxwcuA28gpgKPnoXuJaK37
+GmMkb7+8bxTyfO4yZSkyM+cd+bKiwMa0sHoqr6tnhrcvGzBu9Lp+B9m/LEKmzyjoi45bAd21avr
LsFUam+OOdj2z3RVy+eAjGg/wox0uttYMWwrzJPIjlcF+Sb0gM6muSi3w4v2MoYX8Jlur0g7Ffkq
MQJV30AqI+I6ZvkwnmNlx2Jt6QVXV/6QVX9YCt7OJReJlZUtk6jam28ZXcII7bDlvbJOwCS6W7yt
WpfuF34h9PmdIQmGyqSHZWM/FARnVTNO7LJ1+vml1HiNHNQOSAjK0wiOkIDkxbGN1ijQ0JmdvW9D
khJiIQMGkhOePBJC4GegPSxep6wDpEtT3fbXT88rh2Fwxxc4ATVtPEnl18E5QwcvLKcNa9mpXmxn
2HWjtkHdtdgx73a/D6DpZM7nKNz8omhqavW+KfO/4u/XJDvXLJKQsc1/eNIPVWN+OxaWrZZJJTNk
V2ndhSp0l+EOUYKKZ4W34P3fIU6Tnv5Y4IX5lKA4vswg0zjKtdCKVitF3PKvgisMvdWfDexVDNUZ
NYSqQlc0R5/UdrKHoSjS9zsi1fsQDxZ7E64FrCFuJwLk39JT5uF/ufYNCrV3gX3u8Sf88shNmsCl
ct09XJIHl6t/zwDMFDwaMuC/mGqmQLTClIX4Ztf/PsT6TKNm9DUWKFOM55sosNbKQfvDOMJJrc84
155CDThhjsW3OK7WdXPUlJM02ZGqI5aDGNel2gUt6N/6bxC+4y61l1Iq8TA8xL4hwnkXxuokevhE
ks/4vGwC5e37CCQwLnSLC/YNzuMLbZGFDvUZzwbYxUoDUg0xgkGJZZYUgk690O4bCgxJGBDZKBSQ
72japOqxCTSGb1htsH/GEwL3moYDSId56h7z3zobsjQHMUspxSLwHOyakKUaupt07h1xrIDcyn67
lBrvxlWJndajOfBa3bt/cfHvxGR61XCVO6vwtb/EPiSkf2EpyA7TMUeeWiBuaPV5jRgql4z/1JVQ
u+8lCUq0iv301YvdRQfQBiKH265auNWRHloPkYo5w1C4lO4+N7o4jCp54n5NpSIo7N67jZB38gw7
zUyR0dbSCMno4rUDVLVYI2PQqCzO0pdBoSE/DNxA5QC4KtJTRg1dkEYEiT/aBpQlvLZ0qclCgRDU
VWopSori+VYoS+v2pB+jQS2DjBkb8Iwl22Dtym53KUM8aPpUPMXWNwPvvFBk+7V0HLHGPGCMK+38
1sYbCuiiThHolElunWrSITAyVwqXtG4twH7UgANIZIzoJNA5J+RC0KSr2LlqEC2ITHaD0lKNimOA
X0W2hFjJaRqz4ny1QJxh+xtohzHLfpLq2gfr0WVeOcgYHFzdmAvkQZApEmpVfqHIy6mkaYpOWYO2
MDdaXqPwRoBIWMTu7FPojggM0V+u7XXXi1sR1M8YwmF40IKvJmwRlqGzq9XihC9N4nEQZ4UVLVAP
HsvY4UH83kLXwEDG4KGnfYPaGKIiuQHUAL1AbJbD++rQD1Kt9lPecu5fXRslry+nKzZPmZd1R6nS
bIyTF5N4BuWc+UXdZ6e0HGtiK1ufi0NUThlbDyRouYph5wWnz3g0HANWbbH5FQ+QBSrrmRRyr51L
WM7TzeoqPOmrjG7CZ9NDlQRSNuM1uCetQ6+f7gVy5yUKS7ZSreHU0nG94vEGGGL2IAyRMhYURIxA
uL3C4UOwE3CtqXBZy2vBSYJApMIug/CHdIsFIUMudzJuh49HJA10i2F4RoHYQ9mzCuOBMJdlRi81
SGJUD8E4J05mkp5fKY9sXPrcYffDgmFWqI35pEf4+KvCVK6yg9tgJXM1vbaPVO4O07qdOTrzNY5x
4i6ocFLpeTTioCW3LDhkRurKefw4V0s9KVu541Jzx1Pu9x+MQB1W/2TlDNLH2Zy6sLMRA2cnWC0w
+jfT5c0dnDkneIhye6goyNb2Ju8ewKA9CLlj77j/4UUgcxZgG8PHKCuX2O6FoZLPyF9Ih6tcsRen
0qOS4ekJ2HFQ3vbNr3PVEWDYGB5auEpWBqPCQnhCdjbcJRBU+4pipsAo3i080I3OcCGuBmcL62SM
a1kTDgLnBMbnKuHW65y5kGXtEZBmfKnVCX7POHY5GwuVlPW8EdnF4FwyiMTgGwaDf/ZaJFN3OJuf
3KpCknAeACNt00JJA2bdoh/vTOS56Kj5ec6RDuAT+w4+q0/GTMLPR7Ii1YY/bZ6/ORZZMtdT1PvV
KX4gESTf1IPY/sibyA8E2IhWewYeM2KTde5h3Dk/LVSzzb955ze0qnGCjva/AsF4v3MvskwtxxBk
YENgSa3vI59PMRpM2Cmyhh6qXqK3IJN9NCW+/sAfT+nwFRb4e/JhDo4VaYbfh7wWk41H6sFhbDVv
mIvcR0nQl2ADrabn+xEiBmDSY3AH0wlO6ERE+ajOshtGhsTLBJ9L7C52zLb549Bu83qsOudMkwf5
MTk3iHAo1rgtNBTjmz1kiRzCHXavP0mZE68sFk5O0Iy6NfG/v8P6CNkyyaJXatJkvYdZKYXYhNdw
P3eYlbx4phlD9VhycWrWd30sdMPzxLJE8ZvYaaVwMjzA3pzcTrndjWDIRaI2kRTbmOtt/wRSbUPB
c2sDsV01VRdJognnScbKT5dcMg6IXhsDx4u9Ms7N0czGkynd99u0TE+T61XZdsKgr76GnNvyi/BK
34rXVopkYg8jxstl9XdWqGmFrv8ChZCAElVP0dLeF6734TUSSQbvVkMH3kBakx0HVVlOmAnbzP+/
VKcXngUFSHo1vzPor4B4jJ6q/AgwCt/r+InJyv+dD6VG0fOe0rCPA+4VzcENXaoalsgWGtphdqiL
O7mZMuivBqFcVh6L6nVG520ZIDWSC4oIfAJdtZJ0p9fbXQwnrQMzKxzUR3saWf1dyvAc0ZytEY+j
kGLQ1xB2mVEAqtSHUJsOkzmy389tM1guRJ1J7dfbEhoufidfPAZ3P5AC40teqaetlf4fxAmPg8M3
+/WGQxnKvHnVoB6mE/AYwgOcC4U9hQy7Tifp8x8jJ41CfYQA0wj8vWXg6We7g/bBGgIAEMFoqPEP
VptF9X46lTyrlnFzW7fEzbxvex+4Mv1lecvN9CmG/TcukaID1RW5O8Ol1nmHbPU/s2hmm/1iixVB
/ry3VmQy1aOUPtbPnm6LBqZB/ot8StWJxlg58/ZyOSpOyTYaN/m0b7k11YA4W8d99rSEF8dOVyNv
AvFPnTB9bVeY8EjM7HlP2zj/t3yCWd/I79x3LrKLNpx+frqqYzlSJl4jE/0565XJlEgfmTdzNDhM
M+vSGtGzB9DiUYbySx2nRUavuHvUCA+C12vpxIC5U4M3mpqwUPVOyKzRNRmKDDdPHK2yOi54zetS
dHBwTgcy+hjbixFSon6tI6gZSS7wksY6w3+gQiFvcVNYAKTxipn3mbHTMqW7uCLu4SeOtKyXxeyy
BWJcXzAySQnWtA54HXNom5UIKyYvcowunnBk5HKEXy8u6r9PSaIx/mWx4i9KzLGNFg4/8AzuOUMw
vLjwCisRjvJvynUDP3iPL78uLbIyhZBBx63ksctkPRoHFi07wXIqQ5ePyT0rPSHxblFwfjeHdB2A
+7dnp3eXztUK+d3HSptBie/QuwC9EsqgGoshUZ7NldWXrxOIrwrjyhU0+ByR1VfE85Mz1s66RF/p
QtgtyYArCJ3X+ZsCuigGn9HCL89hmriJ92jb9zNv8f2Os7Nr6fWvIkB19DmVrMEuaqepHKHjUYWo
7uqMn0UQwgMYN08z4URsEL9xgNamrp9GEtWJU9EsvEYMDJEwkXFF6ZN+gR2Nc7QvcE7MonC/FwYQ
cslwURF1D+fHjMEyXLwuM9ZnT7SNZhsMol2MLlgUXiQmfsMu0acCuDC6f9M4nwTVylMuR1GTtbmn
dfqh6fsbD/Iou7OT4GJRmbYTU/aHsoYwN5alpNqAJbZO1w99GbK5fm9O4yH9hoTiAMbCuOD/wg4R
y6Qic5dB6rscOH1FY/Ubsvy5by2s7Uf7SUraAr+v1UUqS9FTurHtZyJNxnheocfEy+efvQbMtPiz
zEA3a+7Qrzk/KvvR6rGIWZZZHIOVuGgKuvkh1ACPMR4v7MsyJTYXOH+l4D86tNrH+J+bprehtbM6
p4ZQLFzsFFN34ZINdKPLGCJn8c7oo0SqbBwbMM60mTR4vIejbaJWoF2eCoJg5noKChcopEnrJitO
ELfm4BkziyqskugqwXOWeZmoEnX8zYCJZmbJjaONDrWgbgWxyf0QksPIrA6CnkEDNypgYR6OwWKQ
9uZnv0jJt7psninR4k3Z/RWn44+Q0Cuz9LAEtItFidVFr6K67h/xPm9GtGr+ek4NdU68gcSJ6G/r
cawLg8smieRkhmXxcXt75+QpQp1F4KV0sySYitsBHWG7mJrbrVJfzr/trQ7R977PHK8/d++3Qi33
wicKtMwf0VqEkjrsYV9z2P9gvTo4siAm5yGsSr4LWmdMT2mIRS2E98HfgnGy+XitvHTS8PVltb3/
vdlIJtOhQVIDHPyM2WDx2Bk4NbyMsgBCXFR67+ewA03wTI2/QqCunCqqD4c7r0tdGV5pAJ3hdVmN
XH+kzMGtGDzwLCiaoW+755mV9pXBEZ36CCB0jGOg8mau2mofOaZgF50fV0qto7/BqORMCgAjDmlG
5MXkRr0lPFn2f7SmYhRkytfzd1T97KMD0hK0ri9kkBe4Ef7lXavGhBKrxXdMiTHDzYPpI36qvNNp
ioTUizJ2bOyg8YNVI5/EyVatd5e0BIgXnRdx1qJ5973cIL4VxuTPaC7LCSR9+b58MvpZYV+jFMo8
57mmVYmUd3HjD7GRJhhTIs4TTMOaklWzbnt5ywcLOwP1NUVCq+2anIks96nnB2Fa+V2EqZYno2Ty
GzSfWmW6waekZ81G6hts8+n58dp4EfDb6q3gQ4WB3LdEMuS6SU97ekVdRGib3ovqCSjFfLrrKct6
cNBGR7WwO9Eus4OFXbF0yOqFNUOPyducfgNYkwBcUZX9mfZ4H9ydEyf02AupUu6Z8q2UxdKjBJqS
04aPg7N9Z5BNNIBzkO3La09q2w6oN84He7hHTELH1XUgVPmi69X+u+Y+lthazYSNRu8KjSC/Py3u
0DeQ5K6EBE3WymOvOr+bfuXOv99n01vWFHvaimcs3AxWpg9X648jag6Dl5aeY8IRSaI6bYBEEqif
AAT1qhysV6exEj0QPmtnB4ON/glmBrqFFGwfG+n5u3BlA6Ntp32zQNCCLgNkc+U1POZ4YssR47CL
YpSNIWYpfrAcmVxH5nrY7jx08FIJ7CKvev4DrFI9C8h+FAjlPr1cqT8cdk7NI6pTw1RhN128zB6g
kTuM6P27xjVd+XEXpfrhsBb3fER7bLhJuColb9yP5egh37bPmDYGsd3O/NCcTJH2S+Sho+mEs3Sv
VUztaHHpjfPUUM1BtoXWVDzQlOy+zEU1dqAvAxmVOoB6LkEv8lFdCovebxD/AIEJLGBe+fMrFvB+
4etXXD3ESzx3htYTOyJbPms5a1zxhW6Gpe++NUf00H3IefNAw3nq0ZZQr5ak3/7Di3k6jb1y9NPq
ruEVUx5c2VfKxk73PB1DmWbdFUJneKuiWk5X183Fh6Ok5SQdnSFtaDrmxeU3elJidKmkQlOMen1J
jzSnqRW6EBs31xzuDmjIftBChgAF8T6uO7f8DChnE4ba1U2upOB86TRBULcTvGKJqN3VSGGC57X7
6TngKXraEsX0cezag5WAfu/YTP89Gb/l7sdaV6/eZYMCSby2nFfFqCWTK5Lh1tMb2GUvUEmYTyDT
tGasLthtOe18BGzN+sqi9dgpoRlEVqC78BihGjpYzkgGUlVPMH0/CgNcldIof1ZG9Qsc0PMinTlt
DrQCmtK6Wa9AJEkWHgaDlxybOvX5p5tFJ3fqwPrYAwSb5GKwPKpknkYw/20xuP3yrKOcT61keBlj
O/Es/lWnhRcL93TWKPYtmKbDSjPYwtkvijvXFD9w0PEDifAjAPEGj2aqX5lNWz6v5JfblOIHFxNp
F+7CodyZ0Hyn6kDj456e6lx7ZFP1CbBQJnIwLFmxty6shCIE3loD+CzUounTRBYmzv5lbD3QQx5L
ikKyBqSKK8MwdyuPhEAzlDrJoZ/3Wx6C+Mje94uosfMDy456PMiNw27UGKcar6XPRGNNqlbDXrrq
e/3SPXnvl6E4IRdHI5isHQ2RDBfZdYJ2wPzCPHbr7gcyryJqAckoOQyNfhYycEJmY2MK79aZgarU
VRScgg1L/Hbwgtw9YVA64MEf1MwTVL0oGbWqjaUxQ31s18yk3L+hlze8QynhGsL9P6ntsltKuW5n
xNbjLt6UodkgM91oO1bwv2zXNxLmeuQkXcdIwrPG0JCZQk8TJXNU6Fljrcyw/65rOtZSrNBtXIKk
l3pr/c+1tYt1jQVXa4pJruCL7R9GiCKmFf4Ge6HuLcl/y1uPBCjysKdHYvWMnBumLfyAwgCHgBNI
aC2a5jKCFUBzAN5dTBbEX2gMlebRclQVn2fAzbGoFf/3FfHc+7rPBc4tl8kOeF6FERcwQUaqLBHj
15f5mSe+K9IVr2yK3zS3Dzy/Wddt7mM0g/ilI5wnUxt74kK23l3dbm8cheztOI+qXKLy4m1FHerv
hQDH1ll/71KrrlzIw7IyhyoZoI1NOGlNV0eJTsOLXTYv0gM3rf7zXk7U/jo/K8cz4e20jDWJHIH3
WC36qjfOjKARFfUMbFxB2qKtpImBwDklTx+prCFJKXD2l68glXwMgGpsUtQNQKK/ptad7pUQ9I7/
qAIPDy0UAWNXxOWpltISCAFP5VoAyEJ3r5ZFhbGPkkR+fnVty+3Y08bayVG6ZQXO/2e03xU4Vdcw
skcANr8O0y/uJwvg3+90VDGd16gAJ7dhJfHfibq/Tvgqc+ZkHsZFSQBnk1pX/0Oz1cURU56Bfyyz
SIKZt3cyfLlRh0Nxp0j6xKKR4nGRBcWT2x4+Fp4VwnELeScGYSQwXFt13zRTF+Ll0L2CdUXiw7xM
TV+mDh6698HkAnKcE3N4/8YqyscWTjdw8R4GzIh916kpNv4EBoqTdZqcuLmTnADg4jPlPe3pD5po
rC4Y1TqvEca9flAsjs+TPcLnNDQwRkdBYBh1ivgmRFY4w5KjSj/jeMFKr3wFezrSilmVQpkAsEWp
RJkeOJWd6CPSjTsepPAUIWOfEnhelq+gZMBR4vTnFYGUngjlW7f24AhbWpbVMZKrJbV8ucso1iWY
TrpAePYpAz4sgTocJFtJ/QAlT6jc7BX7eh9AYJqYSib/y9EhLdd2A8Quh48ZI1p/5XEPAoT2yRYT
9fUAQrykW146V+RRQSWBq1i1p66yqS1+fWB9y60D4JyezIEHpWE2j1kbu7SclFhUnsv6uZbOeT0F
XvJCd/Ydlc+N9ba3XkCZVlNjXWVa9QsSmEEvbXt3vLzUVMj86PEuznUvmpe1pPBYQIFJXMQf8pcQ
9wPK/9w10DsgjRHtvpZlmmcPQhy5VbZ6l88jgb+IggoKEI6nPh8TzC8ehSUbZzIydSIQftZiiiEZ
5z91juHQQs9z7oeR5mYurpamerGWAJCssZTNGyNSJejKfPVyd0X4imdM1lr/mSG+mMn5i01u5IOM
GmPnsXmiFy3h7ipOvJzBEloL0jbSvXOzSqHUlPkrzBPce5XaKYipEjzJQd86v/9ilIh6HS4IYSOk
sr72+JmRx9e1bMr3LcuDG48+GJIDmPMbYGYbtwvwbGGzcM/Wy2piedjiyjs1y6aujCdyw/lGVOAk
HDV1pEajlb07NHM/JFnz4N6rqhQuC2+YauqcRASfHQHOhhOlkmw9QwhFkdLyvJQ6+xkmxzs73m8w
m7Lh96qAcn22UdyYP07qpE3tMgEPlsUy9Gz+8+ft4lSG1RIiyUVmH65aih0pzQhWzYUhjLzhp+pt
d/doTrmu9MtiG1umJQmTtgOjt3vOufWAIDnW4q3/RDHUxiO/a0UvGMSKDuuDv1fAcnwQ8otTvHfd
pfR37x99HMDZF7jLllkxx6DsonG9ZrmTuWUHFWvvbeZzrPL5YJrK6ShCxRIxKNHqPxqYVr3MxC+j
/1BiKUrxPX/s0eBh9NaliQ4u+BndPUWQKpkSqPk0ODiBmmMvVdQMXa5vEzzFysF1OOR2V3bOAZgY
F9YcmnGUHq6g/7pJtfUoa8hefdpzlEoU+t0u6O5XkXvPgaOeK7Z7XqDOvJNW//yh+do8owzQ6Au7
s0Qi2hOR+USYHyWB9zUTsI3GzBbt6P/7JTANMErxmS52A8dIdhACkperHnRcBu4q2P/78IzcZ19L
IxuvnZ/oYm32oZVYuWJEBuQnw7klZJ1GUQfNuOhRk8H18qWSrDAA8kTpRJdkWQ+pEMFKw+6apKV7
3hRgs446akL8F2c6A5OdhGBAqI0ZJB9QxPxBv1jSIN33HyDzVQ7STGG+nISHnPIYrJl4gP4p5VwO
2heZRKSbDzhwBpH7WjatLk/nzOv1lwDM9qR/e3LgRLfK+AGIohE3gQxniOg8kNqspRXQ0kRnPgbc
Wkf8msF5pFiAoGh5w1DdHVvOh5trI1k+lVV+GaQF7TRuTCTyLknnebG5NKHH64kUwZQbUO602aIv
r3Ma5OODIjJIRPJ1py9FjQJiuIq/7UL+P/CJKD3yjEEDqtrm58fuyIFxAl7l9PJkFMSVh+Ii/hL+
jwadZuXQF7UGZJw1+niphphk1k+NcjhybsXFeeZ7Mn5hb9MTzTv5za7eD36CfCQxttK75QGIHljV
ClDYyRYdcIBodgdXj1UYMri82zlp+MjcpqmEsuEgqcOEhcPbjImL0KxK7w88BpALc4H96YmE369J
HsnZ7ytmymm8UZJp0Zj6o8QdfN8orKlYcSTk/3+5AAkDvJmoXGVXD1hwtYZP7IklwTdC7D6XDZbA
YtnPoWdGAuGb9Kf/BVtU8RtDrabq3WCSbCE3kIq8jzR+Z1Z5rxQ8tu0gM/epOzt7O3ZIqAd0qbhV
lu0DKwEK1nss1N6L/FVXT5Jp0aCSfE/17k8uTvAyS/7gbmYkbvLaw21/09+g0vjCE/221B/b/01R
aXUY5UaiMAGgNy4u2xwb3t3bie7TP4mAlTs6qJledYzSIYAizcEW6HCUiBRCbOYsczUEIRuRyvQp
Lmi1mF9fVvw3BTw12b5pyLaQpkh39vIuDWczcawL71CZNH4ytYStJUKldO270sNnl2/NRh6ghGmE
unL3ti0ec3yx/rS+kIAMQNZzfA53V16S7+YBbUXTP1H3NeZMYL/aa4eYhS29Zxrv5j3Mdc8zd5vT
OtPmrSHk/Gw3mk1iWe89ANuXvPIJh4bDYqwW/54U7nkI6vepWLc2N8iKtVThqYYMZjseox6OreyM
WSTQmrjxkMYP/98R33rvRUzJRFpoE9IG28A1eIVuNethXyy6l4b0B4iSCnAtxPbj2Red9woyRiBH
m+6cr2gYHLrrQrNHcghwyEEYeCdusP7vuly73x0zSagpNbYOg0p52FbC5Ehqx3IXNq2FxcJM3auR
a264TKRcH/cbx/0wuVr1XBgYeCC7a2nYRNNChDfvmd0FQ/Crx30qpxe1w79FRWyvE6OCaJjpOjjH
9zFxGx5zuQAv4tpwojvrTePXHPqVjspkuhGCz5biOvrnxtAZPdPJehVd/Z+okHKsZQIqN+n8SXDT
W9vYbNXMoI54zErWPfflqjUGrH3sK77GE/EjY+rr+CFEKZ2I4eJTiWUCm3FldIkV5ivbayMguCm9
MJj+YObXG9vNltTy585Rl89WLVwEvWUVeKniGamdtLOGdPiHimHx3CtuZBexYo6gtwQkqKtFg+QW
shKeJ0ZXqHRYlCu13Zh6xR5AQrb8R/RXu+jroo+F6CFZkkEP5v+zRsB3gPCM2f9Kvzo0Qa0D+k3/
7e0gdBAzMzrcN86MVv+WmMy4F8PmbeKq7UrY1AFdhhNqjkXiu2Fy2fUmzmDc6Ul6717183rrbLkI
OKIQQFkIwk9XApFj+AOz5wdsyY6lfVZspqy+TKhuGm3EbMrbHchAt9Efj8YZh387e0h24tDKM/0s
gTyER9dB3kySzfnMAYdhPazqSoRZm9IOJ9/t+5BCscF5xgbt+OGt7eC37em7PYK4XRX0d/eTD4Dz
WnDvkQdXReJc5Chjha3/I8FJSoVhQ9FhXBx10GzK8PxJyFdGP/9Bvll1ndCi6KLXzRiuMW7CHKun
3QZ88XHWZgsW8r3qXCcBQVYJa4cRMjPyyC9PR7+FMLDwAQR4Uk2ywi72KFyu38bSJg7g3h0+zYp4
MWlc98WK4vEucnivpxB1rpIP8IRRDNd5Poi+kPfA97F/1QFXlyu1QdoB8YBj0ocsrCPa/I8S1het
SARdzVwKPoOES4AO+exKyw/4q4eYzhr5NjWEirRurS7eZjR4YxBIDjn+JTjaYzCa3GkfD/eFV2kk
jNK4K3NsjIAtOBIaRqtu//C+VqBUoTvcyYUFXMFDMQd+jRyX1t3e6LEBDma7rWcXlJSTrbjStAxR
7b0bM4plHwFzUAQaSDpFzRZ6a8kZWgZWXZlJhoSWNTAl1SXEZzk6PXxHey3+5JQpZq2lIqsalkOz
cMiCHoyd50sPfaz+u+9aR5RfbnMPNqAh1BW5GW6ZtfkiGxSsuWBa9GuTuO5lZQuH3MGaSKT3sqKr
fO2AMcN9O9YpMSDLxQ9nF/9MBq46SD1UKSPgkyau71H/RKkj2NMfy6Hp4e+cs8sTs4+qWhw1ACA0
xvLRU6Pwi/u8uYme/qH8HwJrRXmr32PAqqyWS2HKrz4DgSuss3RySsAMPTUndkQdfgxnlgFD5d5M
y8zGHRu6jqNo8H/3wqVzu0wQZECR4Cgi+JsfF8u+gOBsIz9+tT0rW91+HSwWhkdqGIagqwzAuPXY
d7Vy4bgnyGjg56d938O99p5+APZ8Y/5AoVjpvevC0Gm0ANxeJrpnUyp4pu4Ak6aTRThyjWcCeaYz
UwyTQXbx404E0yYAtvQVZl8XBpu5+W7YKko/U6pumoXl3w6DuIMhZG3ebV+OuY+//WEknf2OwtXs
G7rZC1ULaPHn/R3YtZPTkz6aKbOjmFSiP8oMYEGQKhp04f4heREP2j/gabHdClCF7HF3yo4iGBF9
4YB3gpD/TsUrShfD/ZGOr7UDsf4c1fpm9//jIvHTf0gnJnMU0Oy4as1NL1LhlOWpJBixTJOmXyAr
zBvEjxtuakbgF7XhRvzBeZPl6vBxvEnYVUIdNyMs1FOFom+WC3aPIFloGPHHsKPlJkO57jWp7pwo
aemC2cBDmq/adFc+7nctVlamv6cBNz74OfqyXt0c+3jT7F+O2kDxX/+qoGb5mBiSCVBTYmiCSax7
2BLb0+D60F0mggdn+OiEsxmyyRGesXxAeU9S8L8GFbltTA4cp8qmQAXYqpbhqv24/8+1JtDVwi/j
2VyLhidEeBvyQmWCf1lUP1ny2ZgpVVLEB1xfIZC56DaxWY6ZXkG/bqiXgcwe+C3+npCME9Gxkkxf
eNqalwEtVyHRUmJLEodzWgrU8F3zIO9DxfFf5jsZGJTaG6sV2FoGKRTzyXh8ckX7LPSyzk5+ZA/l
livhKMuLh+UjZKwWxiww7Kp+VM93O6Os3glUGqC8Es2zHO3n1qAhoA1ygGPwtKVH0wiiaA+Awk2F
fmahtScaU3oASe7akWMDC1IxuDYx6qyHxuZouaVpDTEDU+4jDycnaQ8Pb/64o8a16FrZ5wKo6ibr
ey9vaQMaXp8iljG28LaiPRj1xcfqawbX7sRT5KhNlEuYBiMd6WgXtXTpUnQbNsJVTMQCEAusGhRf
LPp2SwwXvYrAfVD10Sl7BGyQdWoIeA7BTps8l7QbH0qFdUOnWZb9FZHhfUkjnb7peq7C7uhUdd9M
SmfK784CqIE9EiDIC42afJZWAqhnMxLNZU4oJcmz19C8f9lNJChqTXnXaUAicZqgOxuRLK+33NwX
Qs0XBFRFcvQtuIImzqV250BNfRMePyKRgdA92MvXGIXo+F1DszsjLA0BdiHe4MiivBTX1qN3ODbY
kPFy5zvYCIxTpPzqVuu6YvPCKii9wWwi77ORaV5c9nxVg7gb8jTgFVi2oA08XuJ7oPuKB7a9eRnF
3bx7cgBfhK972mIOfrUoZTRiP9gZlz/RgRugdhhj1NALFJOE95Ua3MNVPYHwn1HjVDvunBhE8Q6v
2LkOJ6iaSyp4RI35vXfEiJsjTQSTD+bPtM/YmsPpT9X7XmDDxlwNf9HedbfQ2GFCgrRcC+y4lQX3
7b63xTkyGMGtjViap/9fgZhI3qOphps297mQDb1g52WndAexFqawCz5vg5RR7riQHe2Q67m2/+xd
l67N2oD6ckmVl25fvQwX2j2kHGofDOWfGDIDr+Mhmc1SJK0DcSD3aIVYYV0v6anKCqdR6sveJ7Ua
BTOa9XJ98HiZ3JPLB72vc9JkT3TgyJJqiabIhhvXIQ+vswO+LoVElKBeQuGDC9cvfmCiioMOJJah
ekWZMLyvFvOOa/iR7hrRuUMZbb+/2wkR/DTohRwVZt/4dNDntKhH3lX70KtcOZgdJahQ8iPqq8l0
iA+rWygIejiCYqPrrWm3cj97WUyGexBt/ROYx4KBEy4EWu/TyTJXo+lFTthsOGHREd8urGRoO7W4
rC/EFZXLwT8Xlc8Sssh9NuC+yE3OWJ/LC2i90XVEkzDDdLpGDXuULeoqy3nf/lDxEfXXaa+oEvXH
v4+stQOOjRTkBtf+31wNymbhO80VktvuoZ4znhscck2VN2jBGkrjWeorIwJnhUG0jnhMbuA+TecY
M7UQ3eKD/ATmDxmurivZgI3OA2XIMeU3lsMYnNTfhcW4ZmyH+n8GvXMVBGpidr96tLKcKRrz8Kob
xqkCfXXIsbYvwy8U/jRgKskUtWs9kLpePaVMFSVso2ZQ38GNvWtlxmuigLIeRfXv4pYi1xiooC3D
Mqoy1fMCr9bFcULsaMhuNeXWdbsts7Zfu9msdjOygEwJh18TfpOyHdQW9nIiYo9NfNKYGY7c+awr
ogehZf3F4H6uOo6Kq9Krs6dpXXe//5SF3PYLnM40/5Fo+pUhwPRU5BvL9FMcoJQgxaIKIs19WUAk
0K8L7gc2idTpKAR3EnEdc4jRvoqPyHH3KU+f8jNHkiT1QQgD5sX0ECuxiCPu1wthwHMv6BZhL0Ah
gmyDeO2qUf8zRaUPgovfYL90481slvH2RoB9y3IhIB+GqGTPaaNyLf3vO3BV85jt2AM4I4AZXQpx
Ch6HnP8haM9wGjWcJhvvuearQjhp4eSoHKXyfOg2mztwwN/I9i0t31h6HjPxITxEpRlW7hN1v2TD
fT9vgm6SrIgEumobOxrURIyABdjl+6F0YVg2HpDLogI/tgNKkxvCfKXnlbYxhLjqBFE3Ku/B31ZS
LlWjdlPP80qvlHUhe+s4ObsvR2/BAg8E9J9r6kHqVn9lbGhJZg0h52HQSdTSiGCE2YOxl+zPDCn3
ifeP36qBTPstPZO5n7ODZAma/Rhgb/xfIndtUp/pcUCv35qNF3I7TOQ9hhcFbmoPBekZTo4Fibxl
cZP9S74IgS5uuxFDleAZN7GhkymhP0sxQeVpbMsRI7iMWyNQlC142GmrfQX/nLZJ5Buo4m1F8ZbI
5GTUptiKoEL7Q1cz6M0l0RTepR19xnISLreS8p9dQaVRrPFHPWgYhiXqNlmvQFQRQXKjAUNBVicc
tSk59PhNn8lDdzJS3imG+Qmujhb+bPxbRhinTm1X8rXHdAcg31OFwSYKAGT9eiKuYbnlmMPj+7bV
3y92JMfo63NvMEBBuMYkzhu2Sq3qHy9FWeidbvl8C2uoY3gaudS0hlWdQgskA2L7oxGl8Cq5T/Sx
pxO6NH+//Q9bx9XwQDvIUbb5ZJmZWbh1a+FRo8Q4cJfMzhPQYo0ZU6vtN/RAOb3K1C0kLsqB+QJK
o8dLvFzlcwQBkV8chrfB72vOQsfWT/1TogEAiYV07hb5Ig/iTj9/VPN+LNCgXmdkLe9S+Q75MBzl
ymXL2zIW0eeKH4y9yOifdgICue9t4NPwVxozO4jVgLn+gm3PCrPVzjcL8IPu27gm8dr6NKVJQp05
jM9BJnT0o8Bi/PKFitRHGoW2JjTzTmq1A6GWKYzzhohXacFepNYW3p/sbyN+jPuySMIn098KYGUD
vHp52usDGXZtEe4qXCy+d6e06DJP1llFxVcX/GDro9s8FEjVa9wXpGsQAtVENSmj2Rm7mR6eJTFK
R2IH82CpglYUNoG3ucutetTTiEpgu5TyqlthdvX1W628FvpBuOhfS9G9pRSXs0GE40a0ew8Xa+Yo
sTsuYIOtNfQ0Va8Qpo3YdEyxxjH85XspJbUq4Ui4PmXYK27Kzx78uLvAqUtb7JhoN6ipLt1ZvHfN
uG3nqKrAWpvtXg3Eg1LqhPtUUKg3Oga5L3E9semcEt7wW5r0N7QSZ6gDhuhx9X51DFb1sQCDK5TK
ifYX3CFhoYCeL67G85RN7WSREWvuPc097ecJEQJK6kX8SxpbIucszl/MehQMNNPjxFHSUG1EFo7G
E+rcgAKLtzGSxjEHMtfmQxDk4w3iilVvnwA4uqViWmEO6GhnL3IdM/vCJyiFFfr5F2k1+w5L/mlN
C7gYSjytQRkFVaidCIZY9IHUqUVHDBimphxizd3sBt/BEMbyHS/E0lFA2y5mrNgTofu5+LkKB+M4
/AhsMkJdmyc0JiiuiOIh9K342vdJwpRnr02wkeXo4z0rbWjS98U1c0oyp+ezGF8suZaAzP2+f9tP
b3RFUeLrtL8vtOyqLQwhLgTaLCUDv8u+OjPurnOQpAacr5u7FRtMl9g6K1IpwITYFuMBPdiYo8/B
1ueSukxl6QK+rmJAGk1L4ecf1ziOKL1y6NdRZXxNeDdchlDY07m04MdX+mWUwCkx3HdbNCwIqfDE
D7xV+1MVwJym7K0YLkELGELP/vKvUxbidRK6etHmf4u1I3uSHBq1zxGBXGQidh4kcDkm7XyeIkQa
AMLXbN6XU/sgscO+F2/6HWaJr26bqG8jVTMDmukNm3Y4Vv+MhLyCUzVrzrZDVAk9rOJnCRhX21qe
+f/vIwI/OfgltnLBy8l5i+KwwHE+8OIHJc1m5Zv/3rhFQtiVYIqxJpw7UxZqjrjxG+XN8nDE1fBN
Hbtb8W+eDTx6BUGKrmO5JABT/tJPX4gM/PzkOrpolTcAAnq54SrGCmuiHF/wSeeFtEHam/knliCC
VkDB79Pokii4dqIOECV0OisBLYxGMlFWUzGeRk7NqzqqvraYmO6z7xBQKLXIK59+4zRKDWOfCDP0
I5CjJ0PcZgC4GNZdytsx2jbLuP7jNCwpROIvm3Fe0HcLrSNiv0N/Z03K5r6Vq1l9KQXE+Dj6+AuU
oXJ6waVOShQUPSvHlk1IrJlJuxKVe84WhfnEngIh/vY1eqOGPGI65ynHkBlF53o6Kw1f/CHcc+uN
gOGRDjZ5pd7RR6Xs+lhsvgnPj/XIuTUlaIG3hIhokfIp81IqhAF2CivbUFMIyz7Tdu8ueuUHah/L
UEC0x4dowkooyI4Dpwp+VkMpjQYzo/Lil8IVjeVr1Don30pvpbmJgacQWr4A1b407s2v51C5pB8/
5hR7kz7ZFcE+VkBE7dnGbE8gRZZGQDCGmMiOsatT9aqojcMCuEldiPSB4JVw/maFGtCh+qEJCTHS
MSW+ivMeka4V20hN7rI8J37S4bTnVYmodT/bzmDxVZ0AqBKe8tqIMUEPKuMwlCohDlW3nKEhMbrC
TTtn02awXIqqlzTuDAorHHaooGjqhH+WX0NJhAvJU7YwCadrmThnJ4bpeM8ZDFG2zWVxjXMJOZ4W
HwzK7+emfSg95kgxTA6SN/KSe1mhsSUiVCcpD+EHX2aYvIkxlQsQovkDyPodXw2FkK9gGLo23A2v
drgNhouq3MLydaKFJ8GKc/CyoAKcaWUoXSUlLVPR6D8hcLJJW66iay9co3SI7Pr6Qrhw3KOUSz8n
FcS18mwzr4TmbeY0+z6CaRQ24O33s9X9CroUlkLusZrAHd0Amd5EF9zE/PVLXRK0kRwOgFMDkibt
/+WwrzB6kZktZ6ZKmplVM8mSg4+Szp47HdheaiG4Us0vPMYG2+RQ1vAFsrAvQQGQEr7qLKQMU40g
1/n/4uaZc/UD5As+fWPGnE7c1MTC09r/cSkKRI+fln4SEzAXJ/hAddfa3AYIcW4fcLP1C7jWgAiw
N0WFPMyDfUAitdMqSLk+HA4YNM1YCd0aM6tZWDb0sTddkgdmTf0ODr4roh4xtSkFF6hFQNhcZeRx
/y8Y2loSe12QOdFRi8yNDlVTImiChiT89unZMlJVc+A46jMBUUCyFDZ0DQb25vQ1z3mn8ovANQuK
89C13vInYA54NNq+Akww5j7CMn3h265A5Ck9MTRvOAkuIqF1Ol6FwjMlXhgSWkzyNc3U8J6tB7S6
9PzARMrXTy0up2ihTdsreSJqWtVBXJBl5mJI5YVSjzO1CZbvQgs1EI+otT15tnbCrDbiHdUIs7sq
UKcKjWZncy/ZfmJkTv4nTMxkGa5jspY9rBWBf2CuQdLSECZqz8NiNumClfSLcGsSOxlFbBhE4LQs
Tv+fba/3EUWClyc4sbOm2MJso/DY7IEJ7fxSSqDXM+ExNgpfr4nf+sk6q7WFi3KJh8ANndhM5I96
qrK2ckgxaXLPMOHqydlJdTVW6JGCsThIJ0WqlJtAWkx8nklVeymHz6yUXnDkHKJQ8nAMc3L8xcch
39vXPbnBYOv0vFjPpg6r262Fo0OgMY+NhEfsAYSjbMyuG7xQdorUiqlUFp7Vt+QuE4w3Ng80WTKA
qxztHxMLpZnIlHMTyqJL1eDTwMxT0riVufdBtXa88BZLM8dnchidQ+f1MgbS9t2QDZG2O3Oxyevy
zclVtVyogz2C7I3/bxLAxuiPhsxx1pQlRq3C5ae1Wlp8ajamJS4gymZd1AhETQFO1phnavRT0pEc
x2mIZpjtvn479NMsmRXLwkcklRPC40324w7ypiJ51r1CmA5OJexgQJXA4QbfGJWq1LiHxxGTxnGb
hIW+qY3XInKNl7TQnjhBO98T/ND7zes/Di7ogQ3cmLWOBBa4JqRDGdbRs9QgZKFTMbk7ma3HtALr
w6CUdHk24iOMvD4QCBNbjbTDwrPFWeStxpeenjvxUAJRzYyGboe/cxTyK5dGbtwYvdD8Kpmzoj0j
VTpsOBcdRv/aNZRVlb43EUYhtFYxkKyvVQisWjPqq8YZcbADKs4Ewv5aquqVDRYruyQtrNo5m129
bKOdWlwI+ZSD32b4np4oprZmSo1R9OEqirM1mP7vapHmXYfH2ZjpdGXcoXGBLJoQRPLllavle/ne
ifOaHbGkQuasAIzRcayXgNGLvgFwZeW4gAS40qCQ3RVe+ZOfmExNPHTBrHK+61hvuAeUpkV58q8h
yF9Xfi2CJ914VhV3ZbMsdG3qPiHINjF7aGINC5x631rljytDfq8X/tLUVhlbu43cqHHUzqe902Rr
lxGpyt/ihNt2eYZ8IsueQLXuATJRikiklGAxZM5JgbZodv/nl48GmBOlY6irUJAQ69uEGdTVbCxo
xBICEalpEHBIyx51S09m1U3RsjPr0I1V1kizS60UzI1rC+MYxO82x1XJ+dVF2h6x2SnZxMMItr1f
wPIHAw5KQ//2RI/bfHVQLyPAcidfdC3yzwAfCSGYZEn6lD/UX56Ol4S0OfItj6DNFBUs4pS3oJZT
90/aGt+vdhC4xUCiOqsKn3DcB4NiEmh4trnaEyg53Hfx9NFdIEVQuv5z8ndCM2PK+DkB4jVe7uyN
8g4rviRHFsIzQw45HpevN0CcJ2+uAID/lzVixlDK6ZjgXU0rSNFXZnRBQFT0yMFRcEKJGUg2s3H2
berz7VQcO7mFd+XwyjPbEmTQ56L6vCCYvYBN1CYg+vUzkFlzJVk6DpY4W2b/xmy/stj1v+kceXkB
qBJI65YxVSYMAdtp/5I2ky8Qnt8PBPXCCp7N5oj3HQ9vbFWIKp/adEUYAvS5krjrLAFoLY0Tnf8/
nNfPIG9oztZXdpCMXvDzLTV7n3R+xgXi0qAH3OgNU5QvpVRpIO20DlxGW8UAwb73KfmvL1QZgM8c
lzeElNUu+QMUjDTPGST8OrodP9o9MA67Rd4t1OtrtUSg/pEpnaqShlVkgg8lwiETAKB/DYqQQp5X
Kz67de5VfIJ4tX60bcDohaIA1T1lcjq1yObZvpNzFafnhvx+OKpqhdCpZgiye1TBv1mcwCNlu1J1
tufJOFqWhhv+RX0uYAkvq7FE+G4Idfd90EdhWCgCuFt31C0wd2Ump5rCdrFhyem6kZdsVXMfBCgp
IchlnVR8Mnv0VQc/RIDQtAf7HQREDk/V6kc881wSO7h2NUq5EqXxb1hexUajGRv5me0xRrjbUF4+
A3PBRK58F9/ced8LieoeWH6jsMc6iwg701yw+UML9Y9X2mj5lcxmiqRBEfaePW9mjcPawgZZT770
DkX0Msif+DZ9q1lTrglKw5SGhlm5v1M1CblElCZ6Sij7hEnjHrZ2Oce/ahAhcT+T1FNAGzqBc4BO
p1rIIqio0FZSTbPafvdtJfrZXNDWF2UGmZnyqKncXe8s7aHJkMTc67+1BcVFUixJQrALq9TnzcJ3
OwBUwf+IK5ZHJ7vjRO9kv4sv7lisHCeng85qRJE6lrp5UA8Dc8SWwtsO6iADVCjdr9vh0JTVAYS4
M3vN54a1clXxQkqWwwbTO0D+tCVHV/ynUILK7TB0uyoyeFJ+c7Sa0iNkMbRvK3XaLBR0frxNvE3D
zy3Rs4kvr3XhN8KAzt4+ytvoavNDt3+jARVPW0Ue3kxvpVvGhD1qp4+cO7bIC5mPdSZc0C7c5Fho
WboasSsjkMj86ec1KhFVa+T8/tb34pXC6xf31E76ajh1XeN+WZqpmYPVMLX6wquQtX7amgf2Vx9G
oRlRT5RifGusC5KPjIo/oqT5hZTQ8jLK5fIbxhVtc4qzWQ2FbzgrnOzVdXNswqW/79h64/dF+Ets
Nw/EKC4OhHqkq2LbPb8hbAZaD1YxoAzqnI2nke1cBZ0wEUEy77JrKGsHKdmYfVhV7s835L1ptnil
nDJHkLzXV4GNBT/dQYDcSO1cMHLlJ2S3b7ZHy57w7U1Lbj72Fm0LrTjCVOQbKe+i78cmt2EIrmmF
9JpMIOVX0cGmytZILfWFHpqqbQrLyCZoMpZj2x3BYIN0ufeppP8hOhDgT+RQSMQVG0TvMlS0UO+A
l3IDh4O6KDZPGI3jrdWNOIhDUHEx7cM0TEx57Jt7QoTvjyj0yDlVmyL8fU2yBApzG1B4LpDuMpLL
IM7L4qGAtZahcbqPf5XLuH9Mbh87Tb6iU6UYz+uwAkJskhP0OLpXF/iAfwyq1t1fCmLJ/TfhjCVg
6Q4gqY3GN6bcqfEZ81o8cjGB4rp49dDvnqFgLlNIRlg5D5i2a83SJF+ZAf9hOMQ+RH2X7YmaVTbr
xYeclKaXvYpMFh/qiXeejduKvDShi3A5NcFeMKRCS5qNGUoPEn6GJbeXO+y1um1Tu93LAoXa0B3z
KxVukAu0k7ZzuH+4sXYf3xDErtt0LtrU9NxbYLVaZyGoqy8fH4bd7NamB8YZPIKxZrzU6T2ClLo3
RIoswehjXl+zBMaPPjvTD8xZqIbYzVwNNItIc4IlK58xD/n7OyEQD4SMvtdvvMtIBTT1fJWYujd4
ACDukPcOlh7plwEyg/XSBOmoCoeGyXTLCgpAMZe1EhVLowLz3TR/ux703KBbXBaNUQYm/rGonOlc
IIiVAhdbrtDw9RvoptLLU9HzDZj+xpNZaHmdhvUDn9i3hx3fF8SF7hivCPAavPJMEPSZhXqSRb01
IA2IEOnHG2tkNyg5kU882zZgVVsCEqjU+nYFtvci+rbDZQLvIel9wPT1cK5bW1NNHcFJqDe2fn3V
3ASOvqm8wruZ4nhIvZrI3n5Q7R84B45ayYTri6XZhc6aG2uxY+jYvzJB+y7vEtHEA+exu/6Xkva9
cIbYpgKj31mDufXDgsl0CaHWAxPIplgO7gMv5gUrU90bLpov4rco6o9lUwN7G/c6+3SthMj+6iYL
IgsgDnZOu1EByIPMt3qupKItxhhxmX/cQakhkV7Jr7m098FvYDkjP94Tgma60ozihu3TzuSGhPrh
dNccI3yfzZ9nnut2yOBB4oZ6S+OKEopQkDgbP3eoS0YGUsvLWy7BrgwuXBbkMEE6VdNwonXsDHvs
m+EFtCb/cPj+s2yyQbnzaWB46RNHY111LLopKeoNZpAt9nO+xzAEJv6CgmDCWQPwdau8dF2ASpxq
UAdBhKgJBgZZyqwSo/ujJuGQiZGi/XvqbxkiDDUZmhH/+yA4OHYTbMOMQ4kCU5KUoOjYoUBMvEz9
kxGLQVICdrHy2yon7OVcF/lRA1TJubsGiMAoxe11tqeOQvjXoP0KA9IxuDTw4tw2OIL0wVKLut7L
/alfCUmn+nsPM63lWlwbo5A4Y1ADe4093ijsDQ7O2AJqrpUGsz1HZqQOCXi8vOXpYWyODRoPVGOR
zGCrPt/AUA0t56yQrsYbk6Yyyvvzy2syR69qprC1GUQM3JjAbOcrQksP9wsN8BsgGn4hXYmaMeuN
PoU3i8W0kNHcftGi7T5qxVmAGeqbcwAEfi6zHyEahnDQBqHqtsaPAyAhcdRsI5otNanNE3/Z9sdX
RDzcFpZ0O2B0O1tPDO2K2Ogn9arF6zDCotA8cMMx0Hdm0RBAEcLst/8mdLkEfEeB/7CMPNsqoBEb
sDU2YpEphemnrnHJFPw/Z7Ruv47rL/y7khbPbMsUXO6D/hI5hHYOxbzjBNYMynqH3CcsD8VjBpLQ
QAJDsermgtFaIih7z6F85/nmTvB8v3Wfxx66qpZQ/8/sdEV8yoWTUY03rBKkaCyHXDBN/9B2GRcZ
8m7Or00tE9qX0LT+eqgRTm2ZJgip1C4HPUgz4HF21nBukzmp+Br1vUnQmROT0wGLNQHdxEzgmr7u
AzHFDZGBz57jXdnLqgnIKNFwQhxMFDGNoWXJ9FqX9qBVLIU2q8Nt8byDKT53mgNERd1ilzz/rPuL
IlAaUsFvhdjpJHCfYaJPbCKZidkrKEXnY+IUGfexI82RVb8tuQnH5/IxG2V4zdjxDGwDYnaD6Gem
X2dLMwHr+bbmBcbX3EqlBiT7P630GEDcFAnQQS0z4mWmi9VssfdLuYFx6pj3POV+cy1Cl/4xZB2L
ZD59hB5h1DeSy8XzHRnm47Cwjaa8C8ND3F+VXN4AUCtrO+8rKPgTNhvdXgjOvSfgRkyXyFl2tJ+V
rIgWC2Um1hh3rN4HnThkf4zIZO3STx1N0V2T8ku5s4SB0/fRDMS2i0fPPrxrhSb2NeaFCfa40vjU
BlP6XFCmvPYkP1+yBL4zSWOmZsYbrXD9ziowhFIX4mMxlD4UxtNyZc5hSZl/04/hL2FvOJUtGZWc
7mypDa75Xa9YxbYuGUPkA+7+FSqdiZsz50M6qRtQljc8fcLlo78BV5aoaINY/4I2xwyi+LKQqztL
UcK8EbRP2ZTP9lgFe6x8u/FGygMJsK2+hjsG90ARh9/+rRV+FM2CkUXTtRFFyWtF6TAL03l63IPs
ZuxFSfBsKjcH46PJ1pnkIiW5UQDDHXReAF2J4ywHphtf8GqhGX4AJ363fNojEEjI8xEYDLAA+g6q
QuvdnU4YxO+yDR0wLjezOuB6764LUaxKLg6vFUBPsLnKhfj2CfnJ9hwciDXsWwDT1PfZaRlvHJkB
mNcO9Q/tZNinj7hNAiCG/0fQ3JbppTKvB1e37+FKqMaOaXfQqO80ivhvY8WetXW94QnnFDBiayM/
cOXfdTvvw1SlC51HZOxXRDGOe381KHOBlCY2P1c5kCBTBOX5/hwO45rO/QlaUwsjRinO6tzlnOxf
hlPZiDjZMGDpP6OSvETdUQ0Npoij/qwqRZ5ugfukzZ484nFxQ5+9t4bg2K7aahISZK77hIy9mP5R
PL4rMMYxj7wlDCDGL9466bQO2G9ko5Lp+vP6o+VsS1+hSfCbHopXdCpBzz1jOy+971wfjAET6xyx
8iY01Cl0NR46YRwk2w==
`protect end_protected
